VERSION 5.7 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
NOWIREEXTENSIONATPIN ON ;
UNITS
  DATABASE MICRONS 1000 ;
  CAPACITANCE PICOFARADS 1000 ;
  CURRENT MILLIAMPS 1000 ;
END UNITS
MANUFACTURINGGRID 0.01 ;
DIVIDERCHAR "/" ;

USEMINSPACING OBS ON ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.01 ;

#------------------------------------------
# ROUTING LAYERS
LAYER ME1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.64 ;
  OFFSET	0 ;
  WIDTH		0.24 ;
  SPACING	0.24 ;
  SPACING   0.28 RANGE 10 1000 ;
  AREA          0.1764 ;
  RESISTANCE	RPERSQ 0.077 ;
  CAPACITANCE	CPERSQDIST 2.593e-05 ;
  EDGECAPACITANCE 9.201e-05 ;
  THICKNESS 0.48 ;
  WIREEXTENSION 0.22 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         0.24 1.0  10.0  20.0 ;
     TABLEENTRIES  2.18 1.48  2.66  2.66 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME1

LAYER VI1
    TYPE CUT ;
    SPACING 0.28 ;
END VI1

LAYER ME2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.64 ;
  OFFSET	0 ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING   0.32 RANGE 10 1000 ;
  AREA          0.1936 ;
  RESISTANCE	RPERSQ 0.062 ;
  CAPACITANCE	CPERSQDIST 1.267e-05 ;
  EDGECAPACITANCE 9.492e-05 ;
  THICKNESS 0.58 ;
  WIREEXTENSION 0.22 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         0.24 1.0  10.0  20.0 ;
     TABLEENTRIES  2.62 1.77  3.25  3.25 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME2

LAYER VI2
    TYPE CUT ;
    SPACING 0.28 ;
END VI2

LAYER ME3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.56  ;
  OFFSET	0  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING   0.32 RANGE 10 1000 ;
  AREA          0.1936 ;
  RESISTANCE	RPERSQ 0.062 ;
  CAPACITANCE	CPERSQDIST 8.163e-06 ;
  EDGECAPACITANCE 9.53e-05 ;
  THICKNESS 0.58 ;
  WIREEXTENSION 0.22 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         0.24 1.0  10.0  20.0 ;
     TABLEENTRIES  2.62 1.77  3.25  3.25 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME3

LAYER VI3
    TYPE CUT ;
    SPACING 0.28 ;
END VI3

LAYER ME4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.64  ;
  OFFSET	0.32  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING   0.32 RANGE 10 1000 ;
  AREA          0.1936 ;
  RESISTANCE	RPERSQ 0.062 ;
  CAPACITANCE	CPERSQDIST 6.021e-06 ;
  EDGECAPACITANCE 9.552e-05 ;
  THICKNESS 0.58 ;
  WIREEXTENSION 0.22 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         0.24 1.0  10.0  20.0 ;
     TABLEENTRIES  2.62 1.77  3.25  3.25 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME4

LAYER VI4
    TYPE CUT ;
    SPACING 0.28 ;
END VI4

LAYER ME5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.56  ;
  OFFSET	0  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING   0.32 RANGE 10 1000 ;
  AREA          0.1936 ;
  RESISTANCE	RPERSQ 0.062 ;
  CAPACITANCE	CPERSQDIST 4.769e-06 ;
  EDGECAPACITANCE 9.557e-05 ;
  THICKNESS 0.58 ;
  WIREEXTENSION 0.22 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         0.24 1.0  10.0  20.0 ;
     TABLEENTRIES  2.62 1.77  3.25  3.25 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME5

LAYER VI5
    TYPE CUT ;
    SPACING 0.28 ;
END VI5

LAYER ME6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		2.2 ;
  OFFSET	0.46 ;
  WIDTH		1.2 ;
  SPACING	1.0 ;
  SPACING   1.5 RANGE 10 1000 ;
  SPACING         0.44 SAMENET ;
  AREA          9.0 ;
  RESISTANCE	RPERSQ 0.02 ;
  CAPACITANCE	CPERSQDIST 3.948e-06 ;
  EDGECAPACITANCE 0.0001047 ;
  THICKNESS 2.06 ;
  WIREEXTENSION 0.54 ;

  DCCURRENTDENSITY AVERAGE
     WIDTH         1.0  10.0  20.0 ;
     TABLEENTRIES  2.96  5.32  5.32 ;

  ANTENNAAREARATIO	400 ;
  ANTENNACUMAREARATIO	 400 ;
  ANTENNAAREAFACTOR	 1 ;
  ANTENNASIDEAREARATIO	 400 ;
  ANTENNACUMSIDEAREARATIO	 400 ;
  ANTENNASIDEAREAFACTOR	 1 ;
END ME6
#------------------------------------------

#------------------------------------------
# DEFINE FOUR DIRECTION DEFAULT VIAS
VIA VIA12_HH DEFAULT
  LAYER ME2 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI1 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME1 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA12_HH
VIA VIA12_HV DEFAULT
  LAYER ME2 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI1 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME1 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA12_HV
VIA VIA12_VH DEFAULT
  LAYER ME2 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI1 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME1 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA12_VH
VIA VIA12_VV DEFAULT
  LAYER ME2 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI1 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME1 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA12_VV
VIA VIA23_HH DEFAULT
  LAYER ME2 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI2 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA23_HH
VIA VIA23_HV DEFAULT
  LAYER ME2 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI2 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA23_HV
VIA VIA23_VH DEFAULT
  LAYER ME2 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI2 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA23_VH
VIA VIA23_VV DEFAULT
  LAYER ME2 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI2 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA23_VV
VIA VIA34_HH DEFAULT
  LAYER ME4 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI3 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA34_HH
VIA VIA34_HV DEFAULT
  LAYER ME4 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI3 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA34_HV
VIA VIA34_VH DEFAULT
  LAYER ME4 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI3 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA34_VH
VIA VIA34_VV DEFAULT
  LAYER ME4 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI3 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME3 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA34_VV
VIA VIA45_HH DEFAULT
  LAYER ME4 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI4 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA45_HH
VIA VIA45_HV DEFAULT
  LAYER ME4 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  LAYER VI4 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA45_HV
VIA VIA45_VH DEFAULT
  LAYER ME4 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI4 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA45_VH
VIA VIA45_VV DEFAULT
  LAYER ME4 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  LAYER VI4 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA45_VV
VIA VIA56_HH DEFAULT
  LAYER ME6 ;
        RECT -0.26 -0.22 0.26 0.22 ;
  LAYER VI5 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA56_HH
VIA VIA56_HV DEFAULT
  LAYER ME6 ;
        RECT -0.26 -0.22 0.26 0.22 ;
  LAYER VI5 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA56_HV
VIA VIA56_VH DEFAULT
  LAYER ME6 ;
        RECT -0.22 -0.26 0.22 0.26 ;
  LAYER VI5 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.22 -0.14 0.22 0.14 ;
  RESISTANCE 6.5 ;
END VIA56_VH
VIA VIA56_VV DEFAULT
  LAYER ME6 ;
        RECT -0.22 -0.26 0.22 0.26 ;
  LAYER VI5 ;
        RECT -0.14 -0.14 0.14 0.14 ;
  LAYER ME5 ;
        RECT -0.14 -0.22 0.14 0.22 ;
  RESISTANCE 6.5 ;
END VIA56_VV
#------------------------------------------

#------------------------------------------
# DEFINE STACK ONLY DEFAULT VIAS
VIA VIA23_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
	 RECT -0.14 -0.48 0.14 0.22 ;
    LAYER VI2 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA23_STACK_HAMMER1
VIA VIA23_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
	 RECT -0.14 -0.22 0.14 0.48 ;
    LAYER VI2 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA23_STACK_HAMMER2
VIA VIA23_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME2 ;
	 RECT -0.14 -0.35 0.14 0.35 ;
    LAYER VI2 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA23_STACK_CROSS
VIA VIA34_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	   RECT -0.14 -0.22 0.14 0.22 ;
    LAYER VI3 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.48 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA34_STACK_HAMMER1
VIA VIA34_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	   RECT -0.14 -0.22 0.14 0.22 ;
    LAYER VI3 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.22 -0.14 0.48 0.14 ;
    RESISTANCE 6.50 ;
END VIA34_STACK_HAMMER2
VIA VIA34_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	   RECT -0.14 -0.22 0.14 0.22 ;
    LAYER VI3 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME3 ;
	   RECT -0.35 -0.14 0.35 0.14 ;
    RESISTANCE 6.50 ;
END VIA34_STACK_CROSS
VIA VIA45_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	 RECT -0.14 -0.48 0.14 0.22 ;
    LAYER VI4 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA45_STACK_HAMMER1
VIA VIA45_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	 RECT -0.14 -0.22 0.14 0.48 ;
    LAYER VI4 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA45_STACK_HAMMER2
VIA VIA45_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME4 ;
	 RECT -0.14 -0.35 0.14 0.35 ;
    LAYER VI4 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.22 -0.14 0.22 0.14 ;
    RESISTANCE 6.50 ;
END VIA45_STACK_CROSS
VIA VIA56_STACK_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER ME6 ;
	   RECT -0.22 -0.26 0.22 0.26 ;
    LAYER VI5 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.44 -0.14 0.26 0.14 ;
    RESISTANCE 6.50 ;
END VIA56_STACK_HAMMER1
VIA VIA56_STACK_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER ME6 ;
	   RECT -0.22 -0.26 0.22 0.26 ;
    LAYER VI5 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.26 -0.14 0.44 0.14 ;
    RESISTANCE 6.50 ;
END VIA56_STACK_HAMMER2
VIA VIA56_STACK_CROSS DEFAULT TOPOFSTACKONLY
    LAYER ME6 ;
	   RECT -0.22 -0.26 0.22 0.26 ;
    LAYER VI5 ;
	   RECT -0.14 -0.14 0.14 0.14 ;
    LAYER ME5 ;
	   RECT -0.35 -0.14 0.35 0.14 ;
    RESISTANCE 6.50 ;
END VIA56_STACK_CROSS

#------------------------------------------
VIA VIA12_HH_2CUT_E DEFAULT 
    LAYER ME1 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_E
VIA VIA12_HH_2CUT_W DEFAULT 
    LAYER ME1 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI1 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_W
VIA VIA12_HH_2CUT_N DEFAULT 
    LAYER ME1 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_N
VIA VIA12_HH_2CUT_S DEFAULT 
    LAYER ME1 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_S
VIA VIA12_HH_2CUT_ALT_E DEFAULT 
    LAYER ME1 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_ALT_E
VIA VIA12_HH_2CUT_ALT_W DEFAULT 
    LAYER ME1 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI1 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_ALT_W
VIA VIA12_HH_2CUT_ALT_N DEFAULT 
    LAYER ME1 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME2 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_ALT_N
VIA VIA12_HH_2CUT_ALT_S DEFAULT 
    LAYER ME1 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    LAYER VI1 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME2 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA12_HH_2CUT_ALT_S
VIA VIA23_HH_MAR_N DEFAULT  TOPOFSTACKONLY
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.220000 0.310000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA23_HH_MAR_N
VIA VIA23_HH_MAR_S DEFAULT  TOPOFSTACKONLY
    LAYER ME2 ; 
	RECT -0.220000 -0.310000 0.220000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA23_HH_MAR_S
VIA VIA23_HH_2CUT_E DEFAULT 
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_E
VIA VIA23_HH_2CUT_W DEFAULT 
    LAYER ME2 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_W
VIA VIA23_HH_2CUT_N DEFAULT 
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_N
VIA VIA23_HH_2CUT_S DEFAULT 
    LAYER ME2 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_S
VIA VIA23_HH_2CUT_ALT_E DEFAULT 
    LAYER ME2 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_ALT_E
VIA VIA23_HH_2CUT_ALT_W DEFAULT 
    LAYER ME2 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI2 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_ALT_W
VIA VIA23_HH_2CUT_ALT_N DEFAULT 
    LAYER ME2 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME3 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_ALT_N
VIA VIA23_HH_2CUT_ALT_S DEFAULT 
    LAYER ME2 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    LAYER VI2 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME3 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA23_HH_2CUT_ALT_S
VIA VIA34_HH_MAR_E DEFAULT  TOPOFSTACKONLY
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.480000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA34_HH_MAR_E
VIA VIA34_HH_MAR_W DEFAULT  TOPOFSTACKONLY
    LAYER ME3 ; 
	RECT -0.480000 -0.140000 0.220000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA34_HH_MAR_W
VIA VIA34_HH_2CUT_E DEFAULT 
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_E
VIA VIA34_HH_2CUT_W DEFAULT 
    LAYER ME3 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_W
VIA VIA34_HH_2CUT_N DEFAULT 
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_N
VIA VIA34_HH_2CUT_S DEFAULT 
    LAYER ME3 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_S
VIA VIA34_HH_2CUT_ALT_E DEFAULT 
    LAYER ME3 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_ALT_E
VIA VIA34_HH_2CUT_ALT_W DEFAULT 
    LAYER ME3 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI3 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_ALT_W
VIA VIA34_HH_2CUT_ALT_N DEFAULT 
    LAYER ME3 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME4 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_ALT_N
VIA VIA34_HH_2CUT_ALT_S DEFAULT 
    LAYER ME3 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    LAYER VI3 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME4 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA34_HH_2CUT_ALT_S
VIA VIA45_HH_MAR_N DEFAULT  TOPOFSTACKONLY
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.220000 0.310000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA45_HH_MAR_N
VIA VIA45_HH_MAR_S DEFAULT  TOPOFSTACKONLY
    LAYER ME4 ; 
	RECT -0.220000 -0.310000 0.220000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 6.500000 ;
END VIA45_HH_MAR_S
VIA VIA45_HH_2CUT_E DEFAULT 
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_E
VIA VIA45_HH_2CUT_W DEFAULT 
    LAYER ME4 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_W
VIA VIA45_HH_2CUT_N DEFAULT 
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_N
VIA VIA45_HH_2CUT_S DEFAULT 
    LAYER ME4 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_S
VIA VIA45_HH_2CUT_ALT_E DEFAULT 
    LAYER ME4 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_ALT_E
VIA VIA45_HH_2CUT_ALT_W DEFAULT 
    LAYER ME4 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI4 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_ALT_W
VIA VIA45_HH_2CUT_ALT_N DEFAULT 
    LAYER ME4 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME5 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_ALT_N
VIA VIA45_HH_2CUT_ALT_S DEFAULT 
    LAYER ME4 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    LAYER VI4 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME5 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA45_HH_2CUT_ALT_S
VIA VIA56_HH_MAR_E DEFAULT  TOPOFSTACKONLY
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.480000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.220000 0.260000 0.220000 ;
    RESISTANCE 6.500000 ;
END VIA56_HH_MAR_E
VIA VIA56_HH_MAR_W DEFAULT  TOPOFSTACKONLY
    LAYER ME5 ; 
	RECT -0.480000 -0.140000 0.220000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.220000 0.260000 0.220000 ;
    RESISTANCE 6.500000 ;
END VIA56_HH_MAR_W
VIA VIA56_HH_2CUT_E DEFAULT 
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.220000 0.820000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_E
VIA VIA56_HH_2CUT_W DEFAULT 
    LAYER ME5 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.820000 -0.220000 0.260000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_W
VIA VIA56_HH_2CUT_N DEFAULT 
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.220000 0.700000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.220000 0.260000 0.780000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_N
VIA VIA56_HH_2CUT_S DEFAULT 
    LAYER ME5 ; 
	RECT -0.220000 -0.700000 0.220000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.780000 0.260000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_S
VIA VIA56_HH_2CUT_ALT_E DEFAULT 
    LAYER ME5 ; 
	RECT -0.220000 -0.140000 0.780000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT 0.420000 -0.140000 0.700000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.260000 -0.220000 0.820000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_ALT_E
VIA VIA56_HH_2CUT_ALT_W DEFAULT 
    LAYER ME5 ; 
	RECT -0.780000 -0.140000 0.220000 0.140000 ;
    LAYER VI5 ; 
	RECT -0.700000 -0.140000 -0.420000 0.140000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.820000 -0.220000 0.260000 0.220000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_ALT_W
VIA VIA56_HH_2CUT_ALT_N DEFAULT 
    LAYER ME5 ; 
	RECT -0.140000 -0.220000 0.140000 0.780000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
	RECT -0.140000 0.420000 0.140000 0.700000 ;
    LAYER ME6 ; 
	RECT -0.220000 -0.260000 0.220000 0.820000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_ALT_N
VIA VIA56_HH_2CUT_ALT_S DEFAULT 
    LAYER ME5 ; 
	RECT -0.140000 -0.780000 0.140000 0.220000 ;
    LAYER VI5 ; 
	RECT -0.140000 -0.700000 0.140000 -0.420000 ;
	RECT -0.140000 -0.140000 0.140000 0.140000 ;
    LAYER ME6 ; 
	RECT -0.220000 -0.820000 0.220000 0.260000 ;
    RESISTANCE 3.250000 ;
END VIA56_HH_2CUT_ALT_S

# END AUTO GENERATED VIAS

VIARULE VIAM1M2A
   LAYER ME1 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.240 TO 0.240 ;
   LAYER ME2 ;
      DIRECTION VERTICAL ;
      WIDTH 0.280 TO 0.280 ;
   VIA VIA12_HH ;
   VIA VIA12_HV ;
   VIA VIA12_VH ;
   VIA VIA12_VV ;
END VIAM1M2A

VIARULE VIAM2M3
   LAYER ME2 ;
      DIRECTION VERTICAL ;
      WIDTH 0.280 TO 0.280 ;
   LAYER ME3 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.280 TO 0.280 ;
   VIA VIA23_HH ;
   VIA VIA23_HV ;
   VIA VIA23_VH ;
   VIA VIA23_VV ;
END VIAM2M3

VIARULE VIAM3M4
   LAYER ME3 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.280 TO 0.280 ;
   LAYER ME4 ;
      DIRECTION VERTICAL ;
      WIDTH 0.280 TO 0.280 ;
   VIA VIA34_HH ;
   VIA VIA34_HV ;
   VIA VIA34_VH ;
   VIA VIA34_VV ;
END VIAM3M4

VIARULE VIAM4M5
   LAYER ME4 ;
      DIRECTION VERTICAL ;
      WIDTH 0.280 TO 0.280 ;
   LAYER ME5 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.280 TO 0.280 ;
   VIA VIA45_HH ;
   VIA VIA45_HV ;
   VIA VIA45_VH ;
   VIA VIA45_VV ;
END VIAM4M5

VIARULE VIAM5M6
   LAYER ME5 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.280 TO 0.280 ;
   LAYER ME6 ;
      DIRECTION VERTICAL ;
      WIDTH 0.440 TO 0.440 ;
   VIA VIA56_HH ;
   VIA VIA56_HV ;
   VIA VIA56_VH ;
   VIA VIA56_VV ;
END VIAM5M6
#------------------------------------------

#------------------------------------------
VIARULE GENM1M2A GENERATE
   LAYER ME1 ;
      WIDTH 0.01 TO 9.99 ;
      ENCLOSURE 0.08 0 ;
   LAYER ME2 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI1 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM1M2A

VIARULE GENM1M2B GENERATE
   LAYER ME1 ;
      WIDTH 10.00 TO 999.0 ;
      ENCLOSURE 0.2 0.2 ;
   LAYER ME2 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI1 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM1M2B

VIARULE GENM2M3A GENERATE
   LAYER ME2 ;
      WIDTH 0.01 TO 9.99 ;
      ENCLOSURE 0.08 0 ;
   LAYER ME3 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI2 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM2M3A

VIARULE GENM2M3B GENERATE
   LAYER ME2 ;
      WIDTH 10.00 TO 999.0 ;
      ENCLOSURE 0.2 0.2 ;
   LAYER ME3 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI2 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM2M3B

VIARULE GENM3M4A GENERATE
   LAYER ME3 ;
      WIDTH 0.01 TO 9.99 ;
      ENCLOSURE 0.08 0 ;
   LAYER ME4 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI3 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM3M4A

VIARULE GENM3M4B GENERATE
   LAYER ME3 ;
      WIDTH 10.00 TO 999.0 ;
      ENCLOSURE 0.2 0.2 ;
   LAYER ME4 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI3 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM3M4B

VIARULE GENM4M5A GENERATE
   LAYER ME4 ;
      WIDTH 0.01 TO 9.99 ;
      ENCLOSURE 0.08 0 ;
   LAYER ME5 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI4 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM4M5A

VIARULE GENM4M5B GENERATE
   LAYER ME4 ;
      WIDTH 10.00 TO 999.0 ;
      ENCLOSURE 0.2 0.2 ;
   LAYER ME5 ;
      ENCLOSURE 0.08 0 ;
   LAYER VI4 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM4M5B

VIARULE GENM5M6A GENERATE
   LAYER ME5 ;
      WIDTH 0.01 TO 9.99 ;
      ENCLOSURE 0.08 0 ;
   LAYER ME6 ;
      ENCLOSURE 0.40 0.40 ;
   LAYER VI5 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM5M6A

VIARULE GENM5M6B GENERATE
   LAYER ME5 ;
      WIDTH 10.00 TO 999.0 ;
      ENCLOSURE 0.2 0.2 ;
   LAYER ME6 ;
      ENCLOSURE 0.40 0.40 ;
   LAYER VI5 ;
      RECT -0.140 -0.140 0.140 0.140 ;
      SPACING 0.560 BY 0.560 ;
END GENM5M6B


SITE CoreSite
  CLASS CORE ;
  SIZE 0.72 BY 5.76 ;
END CoreSite

END LIBRARY
