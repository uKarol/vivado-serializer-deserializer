VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO filterSizeDrawingStyle STRING ;
  MACRO filterSize REAL ;
  MACRO segSnapMode STRING ;
  MACRO snapMode STRING ;
  MACRO ySnapSpacing REAL ;
  MACRO xSnapSpacing REAL ;
  MACRO gridMultiple INTEGER ;
  MACRO gridSpacing REAL ;
  MACRO stopLevel INTEGER ;
  MACRO startLevel INTEGER ;
  MACRO instLabel STRING ;
  MACRO arrayDisplay STRING ;
  MACRO pathCL STRING ;
  MACRO dimmingScope STRING ;
  MACRO dimmingIntensity INTEGER ;
  MACRO instanceDrawingMode STRING ;
  MACRO maxDragFig INTEGER ;
  MACRO maxDragLevel INTEGER ;
  MACRO scrollPercent INTEGER ;
  MACRO lppVisibilityMode STRING ;
END PROPERTYDEFINITIONS

MACRO UCL_AND2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AND2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 3.1 2.02 3.38 2.3 ;
      LAYER ME2 ;
        RECT 3.02 1.94 3.46 2.38 ;
      LAYER ME1 ;
        RECT 3.02 1.94 3.46 2.38 ;
        RECT 3.04 3.56 3.44 4.68 ;
        RECT 3.04 1.08 3.44 1.48 ;
        RECT 3.12 1.08 3.36 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56125 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.170599 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.713217 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.713217 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 6.62576 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 6.62576 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 1.11 1.96 1.51 2.36 ;
        RECT 1.11 1.96 1.44 2.45 ;
        RECT 0.8 2.56 1.23 2.69 ;
        RECT 1.02 2.35 1.11 2.78 ;
        RECT 0.14 2.66 1.02 2.9 ;
        RECT 0.9 2.44 1.35 2.57 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.32 0.44 2.72 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 1.6 1.08 2 1.48 ;
      RECT 1.76 1.08 2 3.1 ;
      RECT 1.4 2.82 1.52 3.28 ;
      RECT 1.28 2.94 2.74 3.1 ;
      RECT 1.52 2.76 1.58 3.16 ;
      RECT 1.24 3.06 2.74 3.1 ;
      RECT 1.58 2.66 2.74 3.1 ;
      RECT 1.12 3.1 1.52 3.28 ;
      RECT 1 3.22 1.4 3.4 ;
      RECT 0.88 3.34 1.28 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_AND2

MACRO UCL_AND2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AND2_2 0 0 ;
  SIZE 4.32 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 3.76 3.56 4.16 5.32 ;
        RECT 0 4.92 4.32 5.32 ;
    END
  END vddd
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.32 0.44 2.72 1.48 ;
        RECT 0 0.44 4.32 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 4.32 5.96 ;
    END
  END vddb
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN1
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 4.32 0.2 ;
    END
  END gndb
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 3.12 1.08 3.36 4.68 ;
        RECT 3.04 1.08 3.44 1.48 ;
        RECT 3.04 3.56 3.44 4.68 ;
        RECT 3.02 1.94 3.46 2.38 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
        RECT 0.9 2.44 1.35 2.57 ;
        RECT 0.14 2.66 1.02 2.9 ;
        RECT 1.02 2.35 1.11 2.78 ;
        RECT 0.8 2.56 1.23 2.69 ;
        RECT 1.11 1.96 1.44 2.45 ;
        RECT 1.11 1.96 1.51 2.36 ;
    END
  END EIN0
  OBS
    LAYER ME1 ;
      RECT 1.6 1.08 2 1.48 ;
      RECT 1.76 1.08 2 3.1 ;
      RECT 1.4 2.82 1.52 3.28 ;
      RECT 1.28 2.94 2.74 3.1 ;
      RECT 1.52 2.76 1.58 3.16 ;
      RECT 1.24 3.06 2.74 3.1 ;
      RECT 1.58 2.66 2.74 3.1 ;
      RECT 1.12 3.1 1.52 3.28 ;
      RECT 1 3.22 1.4 3.4 ;
      RECT 0.88 3.34 1.28 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_AND2_2

MACRO UCL_ANT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_ANT 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.564 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.27 2.88 1.17 3.28 ;
    END
  END A
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
END UCL_ANT

MACRO UCL_AOI21
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AOI21 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.32 0.44 2.72 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.6 3.84 2 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.252 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.7328 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.792 LAYER ME1 ;
    ANTENNADIFFAREA 0.792 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 3.46 0.5 3.74 ;
      LAYER ME2 ;
        RECT 0.14 3.38 0.58 3.82 ;
      LAYER ME1 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.31 2.62 1.12 2.86 ;
        RECT 0.88 1.08 1.12 2.86 ;
        RECT 0.14 3.38 0.58 3.82 ;
        RECT 0.16 4.06 0.56 4.68 ;
        RECT 0.31 2.62 0.55 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2616 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.825758 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.825758 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.181818 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.181818 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.247475 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.247475 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.74 1.94 3.02 ;
      LAYER ME2 ;
        RECT 1.58 2.66 2.02 3.1 ;
      LAYER ME1 ;
        RECT 1.58 2.66 2.02 3.1 ;
        RECT 1.41 2.68 2.02 3.08 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3536 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2576 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.116162 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.116162 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.969697 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.969697 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.247475 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.247475 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 2.02 2.66 2.3 ;
      LAYER ME2 ;
        RECT 2.3 1.94 2.74 2.38 ;
      LAYER ME1 ;
        RECT 2.3 1.94 2.74 2.38 ;
        RECT 2.27 2.38 2.67 2.78 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2056 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8736 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.86532 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.86532 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.676768 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.676768 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 0.14 1.96 0.61 2.36 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN2
  OBS
    LAYER ME1 ;
      RECT 1.04 3.36 2.56 3.6 ;
      RECT 2.32 3.36 2.56 4.68 ;
      RECT 1.04 3.36 1.28 4.68 ;
      RECT 0.88 3.84 1.28 4.68 ;
      RECT 2.32 3.84 2.72 4.68 ;
  END
END UCL_AOI21

MACRO UCL_AOI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AOI22 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7128 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.96 1.24 1.2 4.2 ;
        RECT 0.88 3.38 1.28 4.2 ;
        RECT 0.85 3.38 1.29 3.82 ;
        RECT 1.6 1.08 2 1.48 ;
        RECT 0.96 1.24 2 1.48 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.99 1.96 3.45 2.36 ;
        RECT 3.01 1.94 3.45 2.38 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.29 1.22 2.73 2.02 ;
        RECT 2.21 1.62 2.73 2.02 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
        RECT 0.14 1.96 0.62 2.36 ;
    END
  END EIN2
  PIN EIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.45 2.68 2.01 3.08 ;
        RECT 1.57 2.66 2.01 3.1 ;
    END
  END EIN3
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 2.32 4.32 2.72 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 1.6 3.84 3.44 4.08 ;
      RECT 0.16 3.84 0.56 4.68 ;
      RECT 1.6 3.84 2 4.68 ;
      RECT 0.16 4.44 2 4.68 ;
      RECT 3.04 3.84 3.44 4.68 ;
  END
END UCL_AOI22

MACRO UCL_AOI22_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AOI22_2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.458 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.96 1.24 1.2 4.2 ;
        RECT 0.88 3.38 1.28 4.2 ;
        RECT 0.85 3.38 1.29 3.82 ;
        RECT 1.6 1.08 2 1.48 ;
        RECT 0.96 1.24 2 1.48 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.486 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.99 1.96 3.45 2.36 ;
        RECT 3.01 1.94 3.45 2.38 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.486 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.29 1.22 2.73 2.06 ;
        RECT 2.21 1.66 2.73 2.06 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.486 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
        RECT 0.14 1.96 0.62 2.36 ;
    END
  END EIN2
  PIN EIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.486 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.45 2.68 2.01 3.08 ;
        RECT 1.57 2.66 2.01 3.1 ;
    END
  END EIN3
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 2.32 4.32 2.72 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 1.6 3.84 3.44 4.08 ;
      RECT 0.16 3.56 0.56 4.68 ;
      RECT 1.6 3.56 2 4.68 ;
      RECT 0.16 4.44 2 4.68 ;
      RECT 3.04 3.56 3.44 4.68 ;
  END
END UCL_AOI22_2

MACRO UCL_AON2B
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AON2B 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6908 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.24 1.08 0.48 3.6 ;
        RECT 0.16 1.08 0.56 1.48 ;
        RECT 0.14 2.66 0.58 3.1 ;
        RECT 0.24 3.36 1.2 3.6 ;
        RECT 0.96 3.36 1.2 4.68 ;
        RECT 0.88 3.84 1.28 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.58 1.94 2.02 2.38 ;
        RECT 1.58 1.96 2.23 2.36 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.98 2.68 3.46 3.08 ;
        RECT 3.02 2.66 3.46 3.1 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.73 1.96 1.3 2.36 ;
        RECT 0.86 1.94 1.3 2.38 ;
    END
  END EIN2
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.84 0.56 5.32 ;
        RECT 1.6 3.84 2 5.32 ;
        RECT 3.04 3.84 3.44 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 2.48 1.16 3.44 1.4 ;
      RECT 3.04 1.08 3.44 1.48 ;
      RECT 1.4 2.9 2.72 3.14 ;
      RECT 1.4 2.82 1.77 3.22 ;
      RECT 2.48 1.16 2.72 4.68 ;
      RECT 2.32 3.84 2.72 4.68 ;
  END
END UCL_AON2B

MACRO UCL_AON2B_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_AON2B_2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.24 1.08 0.48 3.1 ;
        RECT 0.16 1.08 0.56 1.48 ;
        RECT 0.14 2.66 0.58 3.1 ;
        RECT 0.14 2.86 1.2 3.1 ;
        RECT 0.96 2.86 1.2 4.68 ;
        RECT 0.88 3.56 1.28 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.58 1.94 2.02 2.38 ;
        RECT 1.58 1.96 2.23 2.36 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.98 2.68 3.46 3.08 ;
        RECT 3.02 2.66 3.46 3.1 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.73 1.96 1.3 2.36 ;
        RECT 0.86 1.94 1.3 2.38 ;
    END
  END EIN2
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 2.48 1.16 3.44 1.4 ;
      RECT 3.04 1.08 3.44 1.48 ;
      RECT 1.45 2.9 2.72 3.14 ;
      RECT 1.45 2.79 1.81 3.19 ;
      RECT 2.48 1.16 2.72 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
  END
END UCL_AON2B_2

MACRO UCL_BUF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF 0 0 ;
  SIZE 4.32 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8304 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9088 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 1.7836 LAYER ME1 ;
    ANTENNADIFFAREA 1.7836 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 3.82 2.02 4.1 2.3 ;
      LAYER ME2 ;
        RECT 3.74 1.94 4.18 2.38 ;
      LAYER ME1 ;
        RECT 2.3 1.94 4.18 2.38 ;
        RECT 3.76 3.56 4.16 4.68 ;
        RECT 3.76 1.08 4.16 1.48 ;
        RECT 3.84 1.08 4.08 4.68 ;
        RECT 2.32 3.56 2.72 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 2.4 1.08 2.64 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 4.32 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 0 4.92 4.32 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 4.32 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 0 0.44 4.32 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 0.96 2.66 2.02 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 3.02 2.66 3.46 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF

MACRO UCL_BUF16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF16 0 0 ;
  SIZE 31.68 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.7232 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 75.0336 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 1.2544 LAYER VI1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 9.58 2.02 9.86 2.3 ;
        RECT 11.02 2.02 11.3 2.3 ;
        RECT 12.46 2.02 12.74 2.3 ;
        RECT 13.9 2.02 14.18 2.3 ;
        RECT 15.34 2.02 15.62 2.3 ;
        RECT 16.78 2.02 17.06 2.3 ;
        RECT 18.22 2.02 18.5 2.3 ;
        RECT 19.66 2.02 19.94 2.3 ;
        RECT 21.1 2.02 21.38 2.3 ;
        RECT 22.54 2.02 22.82 2.3 ;
        RECT 23.98 2.02 24.26 2.3 ;
        RECT 25.42 2.02 25.7 2.3 ;
        RECT 26.86 2.02 27.14 2.3 ;
        RECT 28.3 2.02 28.58 2.3 ;
        RECT 29.74 2.02 30.02 2.3 ;
        RECT 31.18 2.02 31.46 2.3 ;
      LAYER ME2 ;
        RECT 9.5 1.94 31.54 2.38 ;
      LAYER ME1 ;
        RECT 9.5 1.94 31.54 2.38 ;
        RECT 31.12 3.56 31.52 4.68 ;
        RECT 31.12 1.08 31.52 1.48 ;
        RECT 31.2 1.08 31.44 4.68 ;
        RECT 29.68 3.56 30.08 4.68 ;
        RECT 29.68 1.08 30.08 1.48 ;
        RECT 29.76 1.08 30 4.68 ;
        RECT 28.24 3.56 28.64 4.68 ;
        RECT 28.24 1.08 28.64 1.48 ;
        RECT 28.32 1.08 28.56 4.68 ;
        RECT 26.8 3.56 27.2 4.68 ;
        RECT 26.8 1.08 27.2 1.48 ;
        RECT 26.88 1.08 27.12 4.68 ;
        RECT 25.36 3.56 25.76 4.68 ;
        RECT 25.36 1.08 25.76 1.48 ;
        RECT 25.44 1.08 25.68 4.68 ;
        RECT 23.92 3.56 24.32 4.68 ;
        RECT 23.92 1.08 24.32 1.48 ;
        RECT 24 1.08 24.24 4.68 ;
        RECT 22.48 3.56 22.88 4.68 ;
        RECT 22.48 1.08 22.88 1.48 ;
        RECT 22.56 1.08 22.8 4.68 ;
        RECT 21.04 3.56 21.44 4.68 ;
        RECT 21.04 1.08 21.44 1.48 ;
        RECT 21.12 1.08 21.36 4.68 ;
        RECT 19.6 3.56 20 4.68 ;
        RECT 19.6 1.08 20 1.48 ;
        RECT 19.68 1.08 19.92 4.68 ;
        RECT 18.16 3.56 18.56 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.8 1.08 17.04 4.68 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.36 1.08 15.6 4.68 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.48 1.08 12.72 4.68 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 9.52 3.56 9.92 4.68 ;
        RECT 9.52 1.08 9.92 1.48 ;
        RECT 9.6 1.08 9.84 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 31.68 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 7.36 3.56 7.76 5.32 ;
        RECT 8.8 3.56 9.2 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 18.88 3.56 19.28 5.32 ;
        RECT 20.32 3.56 20.72 5.32 ;
        RECT 21.76 3.56 22.16 5.32 ;
        RECT 23.2 3.56 23.6 5.32 ;
        RECT 24.64 3.56 25.04 5.32 ;
        RECT 26.08 3.56 26.48 5.32 ;
        RECT 27.52 3.56 27.92 5.32 ;
        RECT 28.96 3.56 29.36 5.32 ;
        RECT 30.4 3.56 30.8 5.32 ;
        RECT 0 4.92 31.68 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 31.68 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 7.36 0.44 7.76 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 18.88 0.44 19.28 1.48 ;
        RECT 20.32 0.44 20.72 1.48 ;
        RECT 21.76 0.44 22.16 1.48 ;
        RECT 23.2 0.44 23.6 1.48 ;
        RECT 24.64 0.44 25.04 1.48 ;
        RECT 26.08 0.44 26.48 1.48 ;
        RECT 27.52 0.44 27.92 1.48 ;
        RECT 28.96 0.44 29.36 1.48 ;
        RECT 30.4 0.44 30.8 1.48 ;
        RECT 0 0.44 31.68 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 0.96 2.66 2.02 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 2.3 1.94 2.74 2.38 ;
      RECT 2.4 2.66 3.46 3.1 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 4.46 2.66 4.9 3.1 ;
      RECT 5.9 2.66 6.34 3.1 ;
      RECT 7.34 2.66 7.78 3.1 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 5.2 1.08 5.6 1.48 ;
      RECT 6.64 1.08 7.04 1.48 ;
      RECT 8.08 1.08 8.48 1.48 ;
      RECT 3.74 1.94 8.7 2.38 ;
      RECT 8.16 1.94 8.7 3.1 ;
      RECT 8.16 2.66 9.22 3.1 ;
      RECT 3.84 1.08 4.08 4.68 ;
      RECT 5.28 1.08 5.52 4.68 ;
      RECT 6.72 1.08 6.96 4.68 ;
      RECT 8.16 1.08 8.4 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
      RECT 5.2 3.56 5.6 4.68 ;
      RECT 6.64 3.56 7.04 4.68 ;
      RECT 8.08 3.56 8.48 4.68 ;
      RECT 10.22 2.66 10.66 3.1 ;
      RECT 11.66 2.66 12.1 3.1 ;
      RECT 13.1 2.66 13.54 3.1 ;
      RECT 14.54 2.66 14.98 3.1 ;
      RECT 15.98 2.66 16.42 3.1 ;
      RECT 17.42 2.66 17.86 3.1 ;
      RECT 18.86 2.66 19.3 3.1 ;
      RECT 20.3 2.66 20.74 3.1 ;
      RECT 21.74 2.66 22.18 3.1 ;
      RECT 23.18 2.66 23.62 3.1 ;
      RECT 24.62 2.66 25.06 3.1 ;
      RECT 26.06 2.66 26.5 3.1 ;
      RECT 27.5 2.66 27.94 3.1 ;
      RECT 28.94 2.66 29.38 3.1 ;
      RECT 30.38 2.66 30.82 3.1 ;
    LAYER ME2 ;
      RECT 8.16 2.66 30.82 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF16

MACRO UCL_BUF16B
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF16B 0 0 ;
  SIZE 28.8 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 7.36 3.56 7.76 5.32 ;
        RECT 8.8 3.56 9.2 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 18.88 3.56 19.28 5.32 ;
        RECT 20.32 3.56 20.72 5.32 ;
        RECT 21.76 3.56 22.16 5.32 ;
        RECT 23.2 3.56 23.6 5.32 ;
        RECT 24.64 3.56 25.04 5.32 ;
        RECT 26.08 3.56 26.48 5.32 ;
        RECT 27.52 3.56 27.92 5.32 ;
        RECT 0 4.92 28.8 5.32 ;
    END
  END vddd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.7232 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 75.0336 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 1.2544 LAYER VI1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 6.7 2.02 6.98 2.3 ;
        RECT 8.14 2.02 8.42 2.3 ;
        RECT 9.58 2.02 9.86 2.3 ;
        RECT 11.02 2.02 11.3 2.3 ;
        RECT 12.46 2.02 12.74 2.3 ;
        RECT 13.9 2.02 14.18 2.3 ;
        RECT 15.34 2.02 15.62 2.3 ;
        RECT 16.78 2.02 17.06 2.3 ;
        RECT 18.22 2.02 18.5 2.3 ;
        RECT 19.66 2.02 19.94 2.3 ;
        RECT 21.1 2.02 21.38 2.3 ;
        RECT 22.54 2.02 22.82 2.3 ;
        RECT 23.98 2.02 24.26 2.3 ;
        RECT 25.42 2.02 25.7 2.3 ;
        RECT 26.86 2.02 27.14 2.3 ;
        RECT 28.3 2.02 28.58 2.3 ;
      LAYER ME2 ;
        RECT 6.62 1.94 28.66 2.38 ;
      LAYER ME1 ;
        RECT 6.62 1.94 28.66 2.38 ;
        RECT 28.24 3.56 28.64 4.68 ;
        RECT 28.24 1.08 28.64 1.48 ;
        RECT 28.32 1.08 28.56 4.68 ;
        RECT 26.8 3.56 27.2 4.68 ;
        RECT 26.8 1.08 27.2 1.48 ;
        RECT 26.88 1.08 27.12 4.68 ;
        RECT 25.36 3.56 25.76 4.68 ;
        RECT 25.36 1.08 25.76 1.48 ;
        RECT 25.44 1.08 25.68 4.68 ;
        RECT 23.92 3.56 24.32 4.68 ;
        RECT 23.92 1.08 24.32 1.48 ;
        RECT 24 1.08 24.24 4.68 ;
        RECT 22.48 3.56 22.88 4.68 ;
        RECT 22.48 1.08 22.88 1.48 ;
        RECT 22.56 1.08 22.8 4.68 ;
        RECT 21.04 3.56 21.44 4.68 ;
        RECT 21.04 1.08 21.44 1.48 ;
        RECT 21.12 1.08 21.36 4.68 ;
        RECT 19.6 3.56 20 4.68 ;
        RECT 19.6 1.08 20 1.48 ;
        RECT 19.68 1.08 19.92 4.68 ;
        RECT 18.16 3.56 18.56 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.8 1.08 17.04 4.68 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.36 1.08 15.6 4.68 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.48 1.08 12.72 4.68 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 9.52 3.56 9.92 4.68 ;
        RECT 9.52 1.08 9.92 1.48 ;
        RECT 9.6 1.08 9.84 4.68 ;
        RECT 8.08 3.56 8.48 4.68 ;
        RECT 8.08 1.08 8.48 1.48 ;
        RECT 8.16 1.08 8.4 4.68 ;
        RECT 6.64 3.56 7.04 4.68 ;
        RECT 6.64 1.08 7.04 1.48 ;
        RECT 6.72 1.08 6.96 4.68 ;
    END
  END AUS
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 7.36 0.44 7.76 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 18.88 0.44 19.28 1.48 ;
        RECT 20.32 0.44 20.72 1.48 ;
        RECT 21.76 0.44 22.16 1.48 ;
        RECT 23.2 0.44 23.6 1.48 ;
        RECT 24.64 0.44 25.04 1.48 ;
        RECT 26.08 0.44 26.48 1.48 ;
        RECT 27.52 0.44 27.92 1.48 ;
        RECT 0 0.44 28.8 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 28.8 5.96 ;
    END
  END vddb
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7744 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER ME1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.3104 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 28.8 0.2 ;
    END
  END gndb
  OBS
    LAYER ME1 ;
      RECT 1.58 2.66 2.02 3.1 ;
      RECT 3.02 2.66 3.46 3.1 ;
      RECT 4.46 2.66 4.9 3.1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 5.2 1.08 5.6 1.48 ;
      RECT 0.86 1.94 5.82 2.38 ;
      RECT 5.28 1.94 5.82 3.1 ;
      RECT 5.28 2.66 6.34 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 3.84 1.08 4.08 4.68 ;
      RECT 5.28 1.08 5.52 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
      RECT 5.2 3.56 5.6 4.68 ;
      RECT 7.34 2.66 7.78 3.1 ;
      RECT 8.78 2.66 9.22 3.1 ;
      RECT 10.22 2.66 10.66 3.1 ;
      RECT 11.66 2.66 12.1 3.1 ;
      RECT 13.1 2.66 13.54 3.1 ;
      RECT 14.54 2.66 14.98 3.1 ;
      RECT 15.98 2.66 16.42 3.1 ;
      RECT 17.42 2.66 17.86 3.1 ;
      RECT 18.86 2.66 19.3 3.1 ;
      RECT 20.3 2.66 20.74 3.1 ;
      RECT 21.74 2.66 22.18 3.1 ;
      RECT 23.18 2.66 23.62 3.1 ;
      RECT 24.62 2.66 25.06 3.1 ;
      RECT 26.06 2.66 26.5 3.1 ;
      RECT 27.5 2.66 27.94 3.1 ;
    LAYER ME2 ;
      RECT 5.28 2.66 27.94 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF16B

MACRO UCL_BUF4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF4 0 0 ;
  SIZE 7.2 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1008 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3552 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 3.5672 LAYER ME1 ;
    ANTENNADIFFAREA 3.5672 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 6.7 2.02 6.98 2.3 ;
      LAYER ME2 ;
        RECT 6.62 1.94 7.06 2.38 ;
      LAYER ME1 ;
        RECT 2.3 1.94 7.06 2.38 ;
        RECT 6.64 3.56 7.04 4.68 ;
        RECT 6.64 1.08 7.04 1.48 ;
        RECT 6.72 1.08 6.96 4.68 ;
        RECT 5.2 3.56 5.6 4.68 ;
        RECT 5.2 1.08 5.6 1.48 ;
        RECT 5.28 1.08 5.52 4.68 ;
        RECT 3.76 3.56 4.16 4.68 ;
        RECT 3.76 1.08 4.16 1.48 ;
        RECT 3.84 1.08 4.08 4.68 ;
        RECT 2.32 3.56 2.72 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 2.4 1.08 2.64 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 7.2 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 0 4.92 7.2 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 7.2 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 0 0.44 7.2 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 0.96 2.66 2.02 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 3.02 2.66 3.46 3.1 ;
      RECT 4.46 2.66 4.9 3.1 ;
      RECT 5.9 2.66 6.34 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF4

MACRO UCL_BUF8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF8 0 0 ;
  SIZE 18.72 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6416 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 37.248 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.6272 LAYER VI1 ;
    ANTENNADIFFAREA 7.1344 LAYER ME1 ;
    ANTENNADIFFAREA 7.1344 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 8.14 2.02 8.42 2.3 ;
        RECT 9.58 2.02 9.86 2.3 ;
        RECT 11.02 2.02 11.3 2.3 ;
        RECT 12.46 2.02 12.74 2.3 ;
        RECT 13.9 2.02 14.18 2.3 ;
        RECT 15.34 2.02 15.62 2.3 ;
        RECT 16.78 2.02 17.06 2.3 ;
        RECT 18.22 2.02 18.5 2.3 ;
      LAYER ME2 ;
        RECT 8.06 1.94 18.58 2.38 ;
      LAYER ME1 ;
        RECT 8.06 1.94 18.58 2.38 ;
        RECT 18.16 3.56 18.56 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.8 1.08 17.04 4.68 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.36 1.08 15.6 4.68 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.48 1.08 12.72 4.68 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 9.52 3.56 9.92 4.68 ;
        RECT 9.52 1.08 9.92 1.48 ;
        RECT 9.6 1.08 9.84 4.68 ;
        RECT 8.08 3.56 8.48 4.68 ;
        RECT 8.08 1.08 8.48 1.48 ;
        RECT 8.16 1.08 8.4 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 18.72 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 7.36 3.56 7.76 5.32 ;
        RECT 8.8 3.56 9.2 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 0 4.92 18.72 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 18.72 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 7.36 0.44 7.76 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 0 0.44 18.72 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 0.96 2.66 2.02 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 2.3 1.94 2.74 2.38 ;
      RECT 2.4 2.66 3.46 3.1 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 4.46 2.66 4.9 3.1 ;
      RECT 5.9 2.66 6.34 3.1 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 5.2 1.08 5.6 1.48 ;
      RECT 6.64 1.08 7.04 1.48 ;
      RECT 3.74 1.94 7.26 2.38 ;
      RECT 6.72 1.94 7.26 3.1 ;
      RECT 6.72 2.66 7.78 3.1 ;
      RECT 3.84 1.08 4.08 4.68 ;
      RECT 5.28 1.08 5.52 4.68 ;
      RECT 6.72 1.08 6.96 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
      RECT 5.2 3.56 5.6 4.68 ;
      RECT 6.64 3.56 7.04 4.68 ;
      RECT 8.78 2.66 9.22 3.1 ;
      RECT 10.22 2.66 10.66 3.1 ;
      RECT 11.66 2.66 12.1 3.1 ;
      RECT 13.1 2.66 13.54 3.1 ;
      RECT 14.54 2.66 14.98 3.1 ;
      RECT 15.98 2.66 16.42 3.1 ;
      RECT 17.42 2.66 17.86 3.1 ;
    LAYER ME2 ;
      RECT 6.72 2.66 17.86 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF8

MACRO UCL_BUF8_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_BUF8_2 0 0 ;
  SIZE 15.84 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6416 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 37.248 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.6272 LAYER VI1 ;
    ANTENNADIFFAREA 7.1344 LAYER ME1 ;
    ANTENNADIFFAREA 7.1344 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 5.26 2.02 5.54 2.3 ;
        RECT 6.7 2.02 6.98 2.3 ;
        RECT 8.14 2.02 8.42 2.3 ;
        RECT 9.58 2.02 9.86 2.3 ;
        RECT 11.02 2.02 11.3 2.3 ;
        RECT 12.46 2.02 12.74 2.3 ;
        RECT 13.9 2.02 14.18 2.3 ;
        RECT 15.34 2.02 15.62 2.3 ;
      LAYER ME2 ;
        RECT 5.18 1.94 15.7 2.38 ;
      LAYER ME1 ;
        RECT 5.18 1.94 15.7 2.38 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.36 1.08 15.6 4.68 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.48 1.08 12.72 4.68 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 9.52 3.56 9.92 4.68 ;
        RECT 9.52 1.08 9.92 1.48 ;
        RECT 9.6 1.08 9.84 4.68 ;
        RECT 8.08 3.56 8.48 4.68 ;
        RECT 8.08 1.08 8.48 1.48 ;
        RECT 8.16 1.08 8.4 4.68 ;
        RECT 6.64 3.56 7.04 4.68 ;
        RECT 6.64 1.08 7.04 1.48 ;
        RECT 6.72 1.08 6.96 4.68 ;
        RECT 5.2 3.56 5.6 4.68 ;
        RECT 5.2 1.08 5.6 1.48 ;
        RECT 5.28 1.08 5.52 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5808 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5344 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9828 LAYER ME1 ;
      ANTENNAGATEAREA 0.9828 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.079772 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.079772 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 15.84 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 7.36 3.56 7.76 5.32 ;
        RECT 8.8 3.56 9.2 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 0 4.92 15.84 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 15.84 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 7.36 0.44 7.76 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 0 0.44 15.84 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 1.58 2.66 2.02 3.1 ;
      RECT 3.02 2.66 3.46 3.1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 0.86 1.94 4.38 2.38 ;
      RECT 3.84 1.94 4.38 3.1 ;
      RECT 3.84 2.66 4.9 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 3.84 1.08 4.08 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
      RECT 5.9 2.66 6.34 3.1 ;
      RECT 7.34 2.66 7.78 3.1 ;
      RECT 8.78 2.66 9.22 3.1 ;
      RECT 10.22 2.66 10.66 3.1 ;
      RECT 11.66 2.66 12.1 3.1 ;
      RECT 13.1 2.66 13.54 3.1 ;
      RECT 14.54 2.66 14.98 3.1 ;
    LAYER ME2 ;
      RECT 3.84 2.66 14.98 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_BUF8_2

MACRO UCL_CAP5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CAP5 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.6 4.64 2 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.2 0.44 1.6 4.18 ;
        RECT 2 0.44 2.4 4.18 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_CAP5

MACRO UCL_CAP6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CAP6 0 0 ;
  SIZE 4.32 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 4.32 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.71 4.42 2.61 5.32 ;
        RECT 0 4.92 4.32 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 4.32 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.2 0.44 1.6 4.18 ;
        RECT 2.72 0.44 3.12 4.18 ;
        RECT 0 0.44 4.32 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_CAP6

MACRO UCL_CAP7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CAP7 0 0 ;
  SIZE 5.04 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 5.04 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 2.07 4.42 2.97 5.32 ;
        RECT 0 4.92 5.04 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 5.04 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.2 0.44 1.6 4.18 ;
        RECT 3.44 0.44 3.84 4.18 ;
        RECT 0 0.44 5.04 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_CAP7

MACRO UCL_CAP8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CAP8 0 0 ;
  SIZE 5.76 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 5.76 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 2.43 4.42 3.33 5.32 ;
        RECT 0 4.92 5.76 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 5.76 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.2 0.44 1.6 4.18 ;
        RECT 4.16 0.44 4.56 4.18 ;
        RECT 0 0.44 5.76 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_CAP8

MACRO UCL_CAP9
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CAP9 0 0 ;
  SIZE 6.48 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 6.48 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 2.79 4.42 3.69 5.32 ;
        RECT 0 4.92 6.48 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 6.48 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.2 0.44 1.6 4.18 ;
        RECT 4.88 0.44 5.28 4.18 ;
        RECT 0 0.44 6.48 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_CAP9

MACRO UCL_CGI2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_CGI2 0 0 ;
  SIZE 4.32 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2056 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8736 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.313797 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.313797 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 1.333333 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 1.333333 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.82 2.02 4.1 2.3 ;
      LAYER ME2 ;
        RECT 3.74 1.94 4.18 2.38 ;
      LAYER ME1 ;
        RECT 3.74 1.94 4.18 2.38 ;
        RECT 3.71 1.96 4.18 2.36 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3776 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2864 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.2376 LAYER ME1 ;
    ANTENNADIFFAREA 0.9828 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 3.86 2.66 4.14 ;
        RECT 2.38 1.3 2.66 1.58 ;
      LAYER ME2 ;
        RECT 2.3 3.78 2.74 4.22 ;
        RECT 2.3 1.22 2.74 1.66 ;
        RECT 2.38 1.22 2.66 4.22 ;
      LAYER ME1 ;
        RECT 2.3 1.22 2.74 1.66 ;
        RECT 2.32 1.08 2.72 1.66 ;
        RECT 2.3 3.78 2.74 4.22 ;
        RECT 2.32 3.78 2.72 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0464 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.436508 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.436508 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 1.59707 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 1.59707 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.68 0.5 2.96 ;
      LAYER ME2 ;
        RECT 0.14 2.6 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.6 0.79 3.04 ;
    END
  END EIN0
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2616 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.798535 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.798535 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.1 2.68 3.38 2.96 ;
      LAYER ME2 ;
        RECT 3.02 2.6 3.46 3.1 ;
      LAYER ME1 ;
        RECT 2.85 2.64 3.46 3.04 ;
        RECT 3.02 2.6 3.46 3.04 ;
    END
  END EIN2
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 4.32 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.78 1.28 5.32 ;
        RECT 3.76 3.56 4.16 5.32 ;
        RECT 0 4.92 4.32 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 4.32 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 3.76 0.44 4.16 1.48 ;
        RECT 0 0.44 4.32 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.24 3.28 3.36 3.52 ;
      RECT 3.04 3.28 3.36 4.68 ;
      RECT 0.24 3.28 0.48 4.68 ;
      RECT 0.16 3.78 0.56 4.68 ;
      RECT 3.04 3.56 3.44 4.68 ;
      RECT 0.16 1.08 0.56 1.48 ;
      RECT 3.04 1.08 3.44 1.48 ;
      RECT 0.24 1.08 0.48 2.14 ;
      RECT 3.16 1.08 3.4 2.14 ;
      RECT 0.24 1.9 3.4 2.14 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_CGI2

MACRO UCL_DELAY
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DELAY 0 0 ;
  SIZE 7.2 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 7.2 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 4.28 0.56 5.32 ;
        RECT 2.06 4.28 2.46 5.32 ;
        RECT 3.96 4.28 4.36 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 0 4.92 7.2 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 7.2 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.06 0.44 2.46 1.48 ;
        RECT 3.96 0.44 4.36 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 0 0.44 7.2 0.84 ;
    END
  END gndd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 6.72 1.08 6.96 4.68 ;
        RECT 6.64 1.08 7.04 1.48 ;
        RECT 6.64 3.56 7.04 4.68 ;
        RECT 6.62 1.94 7.06 2.38 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.34 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  OBS
    LAYER ME1 ;
      RECT 1.34 2.76 2.46 3 ;
      RECT 2.06 2.68 2.46 3.08 ;
      RECT 1.34 1.08 1.74 4.68 ;
      RECT 3.24 2.76 4.36 3 ;
      RECT 3.96 2.68 4.36 3.08 ;
      RECT 3.24 1.08 3.64 4.68 ;
      RECT 5.14 2.76 6.34 3 ;
      RECT 5.9 2.66 6.34 3.1 ;
      RECT 5.14 1.08 5.54 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_DELAY

MACRO UCL_DFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF 0 0 ;
  SIZE 14.4 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 14.4 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.5 0.44 0.9 1.48 ;
        RECT 2.86 0.44 3.26 1.48 ;
        RECT 5.78 0.44 6.18 1.48 ;
        RECT 9.06 0.44 9.46 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 0 0.44 14.4 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 14.4 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.22 3.56 1.62 5.32 ;
        RECT 3.58 3.56 3.98 5.32 ;
        RECT 5.78 3.56 6.18 5.32 ;
        RECT 8.4 3.59 8.8 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 0 4.92 14.4 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 7.42 2.02 7.7 2.3 ;
      LAYER ME2 ;
        RECT 7.34 1.94 7.78 2.38 ;
      LAYER ME1 ;
        RECT 7.34 1.94 7.78 2.38 ;
        RECT 7.07 1.66 7.64 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9322 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025199 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 2.845543 LAYER ME1 ;
      ANTENNAMAXAREACAR 2.845543 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 9.234429 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 9.234429 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.49 2.8 1.89 3.2 ;
        RECT 1.49 2.34 1.73 3.2 ;
        RECT 1.25 2.22 1.61 2.44 ;
        RECT 1.13 2.1 1.49 2.32 ;
        RECT 1.37 2.34 1.73 2.56 ;
        RECT 0.14 1.98 1.37 2.14 ;
        RECT 0.14 1.86 1.25 2.14 ;
        RECT 0.14 1.74 1.13 2.14 ;
        RECT 1.07 2.1 1.49 2.2 ;
        RECT 0.14 1.74 0.73 2.38 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 12.46 2.02 12.74 2.3 ;
      LAYER ME2 ;
        RECT 12.38 1.94 12.82 2.38 ;
      LAYER ME1 ;
        RECT 12.38 1.94 12.82 2.38 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.51 1.08 12.75 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 13.9 2.74 14.18 3.02 ;
      LAYER ME2 ;
        RECT 13.82 2.66 14.26 3.1 ;
      LAYER ME1 ;
        RECT 13.82 2.66 14.26 3.1 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 1.68 1.08 2.08 1.48 ;
      RECT 1.84 1.08 2.08 1.84 ;
      RECT 1.96 1.74 3.75 1.96 ;
      RECT 2.08 1.74 3.75 1.98 ;
      RECT 2.08 1.62 2.18 2.06 ;
      RECT 3.35 1.74 3.75 2.14 ;
      RECT 2.18 2.72 2.54 2.85 ;
      RECT 2.18 1.72 2.2 2.85 ;
      RECT 2.2 1.74 2.42 2.97 ;
      RECT 2.32 2.84 2.64 3.05 ;
      RECT 2.4 2.84 2.64 4.68 ;
      RECT 2.4 3.56 2.8 4.68 ;
      RECT 3.58 1.08 3.98 1.48 ;
      RECT 3.58 1.31 4.51 1.48 ;
      RECT 3.58 1.24 4.39 1.48 ;
      RECT 4.2 1.43 4.63 1.6 ;
      RECT 4.32 1.43 4.63 1.67 ;
      RECT 4.39 1.87 4.87 2.27 ;
      RECT 2.67 2.22 3.07 2.62 ;
      RECT 2.67 2.38 4.63 2.62 ;
      RECT 4.39 1.43 4.63 4.68 ;
      RECT 4.3 3.56 4.7 4.68 ;
      RECT 5.59 2.83 6 3.2 ;
      RECT 5.59 3.04 6.62 3.2 ;
      RECT 5.59 2.96 6.5 3.2 ;
      RECT 6.32 3.16 6.74 3.3 ;
      RECT 6.42 3.28 6.86 3.38 ;
      RECT 6.5 3.28 6.86 4.68 ;
      RECT 6.5 3.4 6.9 4.68 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.46 1.68 6.74 1.84 ;
      RECT 6.5 1.08 6.74 1.84 ;
      RECT 5.59 1.72 6.69 1.96 ;
      RECT 5.59 1.72 5.99 2.11 ;
      RECT 5.06 1.08 5.46 1.48 ;
      RECT 5.11 2.35 7.09 2.59 ;
      RECT 6.69 2.35 7.09 2.87 ;
      RECT 6.69 2.63 9.76 2.87 ;
      RECT 4.87 2.6 5.35 3 ;
      RECT 9.36 2.63 9.76 3.09 ;
      RECT 5.11 1.08 5.35 4.68 ;
      RECT 5.06 3.56 5.46 4.68 ;
      RECT 7.88 1.08 8.28 1.48 ;
      RECT 10.24 1.08 10.64 1.48 ;
      RECT 8.11 1.08 8.28 1.6 ;
      RECT 8.23 1.54 8.59 1.65 ;
      RECT 8.28 1.61 8.7 1.77 ;
      RECT 9.69 1.59 10.24 1.96 ;
      RECT 9.57 1.6 10.24 1.96 ;
      RECT 8.28 1.3 8.4 1.77 ;
      RECT 8.4 1.42 8.52 1.89 ;
      RECT 9.7 1.24 10.24 1.96 ;
      RECT 8.52 1.72 10.24 1.96 ;
      RECT 10 2.15 10.94 2.55 ;
      RECT 9.05 3.13 9.17 3.8 ;
      RECT 7.74 3.11 9.05 3.35 ;
      RECT 7.62 3.21 7.74 3.67 ;
      RECT 7.51 3.33 7.94 3.45 ;
      RECT 8.93 3.25 9.29 3.45 ;
      RECT 9.03 3.25 9.29 3.47 ;
      RECT 7.39 3.44 7.84 3.55 ;
      RECT 7.39 3.44 7.74 3.67 ;
      RECT 9.05 3.25 9.29 3.8 ;
      RECT 10 1.24 10.24 3.8 ;
      RECT 9.05 3.56 10.24 3.8 ;
      RECT 7.22 3.56 7.62 4.68 ;
      RECT 9.58 3.56 9.98 4.68 ;
      RECT 10.96 1.08 11.36 1.48 ;
      RECT 11.12 1.08 11.36 1.85 ;
      RECT 11.18 2.15 11.8 2.55 ;
      RECT 11.18 1.66 11.43 3.5 ;
      RECT 11.11 3.34 11.36 4.68 ;
      RECT 10.96 3.56 11.36 4.68 ;
  END
END UCL_DFF

MACRO UCL_DFF_LP
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_LP 0 0 ;
  SIZE 14.4 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 14.4 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.5 0.44 0.9 1.48 ;
        RECT 2.85 0.44 3.25 1.08 ;
        RECT 2.86 1.08 3.26 1.48 ;
        RECT 5.78 0.44 6.18 1.48 ;
        RECT 9.06 0.44 9.46 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 0 0.44 14.4 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 14.4 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.22 4.28 1.62 5.32 ;
        RECT 3.58 4.28 3.98 5.32 ;
        RECT 5.78 3.84 6.18 5.32 ;
        RECT 8.4 4.28 8.8 5.32 ;
        RECT 11.68 4.28 12.08 5.32 ;
        RECT 13.12 4.28 13.52 5.32 ;
        RECT 0 4.92 14.4 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 7.42 2.02 7.7 2.3 ;
      LAYER ME2 ;
        RECT 7.34 1.94 7.78 2.38 ;
      LAYER ME1 ;
        RECT 7.34 1.94 7.78 2.38 ;
        RECT 7.07 1.66 7.64 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9322 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025199 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME2 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME1 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.49 2.8 1.89 3.2 ;
        RECT 1.49 2.34 1.73 3.2 ;
        RECT 1.25 2.22 1.61 2.44 ;
        RECT 1.13 2.1 1.49 2.32 ;
        RECT 1.37 2.34 1.73 2.56 ;
        RECT 0.14 1.98 1.37 2.14 ;
        RECT 0.14 1.86 1.25 2.14 ;
        RECT 0.14 1.74 1.13 2.14 ;
        RECT 1.07 2.1 1.49 2.2 ;
        RECT 0.14 1.74 0.73 2.38 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 12.46 2.02 12.74 2.3 ;
      LAYER ME2 ;
        RECT 12.38 1.94 12.82 2.38 ;
      LAYER ME1 ;
        RECT 12.38 1.94 12.82 2.38 ;
        RECT 12.4 4.28 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.51 1.08 12.75 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 13.9 2.74 14.18 3.02 ;
      LAYER ME2 ;
        RECT 13.82 2.66 14.26 3.1 ;
      LAYER ME1 ;
        RECT 13.82 2.66 14.26 3.1 ;
        RECT 13.84 4.28 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 1.68 1.08 2.08 1.48 ;
      RECT 1.84 1.08 2.08 1.84 ;
      RECT 1.96 1.74 3.75 1.96 ;
      RECT 2.08 1.74 3.75 1.98 ;
      RECT 2.08 1.62 2.18 2.06 ;
      RECT 3.35 1.74 3.75 2.14 ;
      RECT 2.18 2.72 2.54 2.85 ;
      RECT 2.18 1.72 2.2 2.85 ;
      RECT 2.2 1.74 2.42 2.97 ;
      RECT 2.32 2.84 2.64 3.05 ;
      RECT 2.4 2.84 2.64 4.68 ;
      RECT 2.4 4.28 2.8 4.68 ;
      RECT 3.58 1.08 3.98 1.48 ;
      RECT 3.58 1.31 4.51 1.48 ;
      RECT 3.58 1.24 4.39 1.48 ;
      RECT 4.2 1.43 4.63 1.6 ;
      RECT 4.32 1.43 4.63 1.67 ;
      RECT 4.39 1.87 4.87 2.27 ;
      RECT 2.67 2.22 3.07 2.62 ;
      RECT 2.67 2.38 4.63 2.62 ;
      RECT 4.39 1.43 4.63 4.68 ;
      RECT 4.3 4.28 4.7 4.68 ;
      RECT 5.59 2.83 6 3.2 ;
      RECT 5.59 3.04 6.62 3.2 ;
      RECT 5.59 2.96 6.5 3.2 ;
      RECT 6.32 3.16 6.74 3.3 ;
      RECT 6.42 3.28 6.86 3.38 ;
      RECT 6.5 3.28 6.86 4.68 ;
      RECT 6.5 3.4 6.9 4.68 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.46 1.68 6.74 1.84 ;
      RECT 6.5 1.08 6.74 1.84 ;
      RECT 5.59 1.72 6.69 1.96 ;
      RECT 5.59 1.72 5.99 2.11 ;
      RECT 5.06 1.08 5.46 1.48 ;
      RECT 5.11 2.35 7.09 2.59 ;
      RECT 6.69 2.35 7.09 2.87 ;
      RECT 6.69 2.63 9.76 2.87 ;
      RECT 4.87 2.6 5.35 3 ;
      RECT 9.36 2.63 9.76 3.09 ;
      RECT 5.11 1.08 5.35 4.68 ;
      RECT 5.06 3.84 5.46 4.68 ;
      RECT 7.88 1.08 8.28 1.48 ;
      RECT 10.24 1.08 10.64 1.48 ;
      RECT 8.11 1.08 8.28 1.6 ;
      RECT 8.23 1.54 8.59 1.65 ;
      RECT 8.28 1.61 8.7 1.77 ;
      RECT 9.69 1.59 10.24 1.96 ;
      RECT 9.57 1.6 10.24 1.96 ;
      RECT 8.28 1.3 8.4 1.77 ;
      RECT 8.4 1.42 8.52 1.89 ;
      RECT 9.7 1.24 10.24 1.96 ;
      RECT 8.52 1.72 10.24 1.96 ;
      RECT 10 2.15 10.94 2.55 ;
      RECT 9.05 3.13 9.17 3.8 ;
      RECT 7.74 3.11 9.05 3.35 ;
      RECT 7.62 3.21 7.74 3.67 ;
      RECT 7.51 3.33 7.94 3.45 ;
      RECT 8.93 3.25 9.29 3.45 ;
      RECT 9.03 3.25 9.29 3.47 ;
      RECT 7.39 3.44 7.84 3.55 ;
      RECT 7.39 3.44 7.74 3.67 ;
      RECT 9.05 3.25 9.29 3.8 ;
      RECT 10 1.24 10.24 3.8 ;
      RECT 9.05 3.56 10.24 3.8 ;
      RECT 7.22 3.56 7.62 4.68 ;
      RECT 9.58 3.56 9.98 4.68 ;
      RECT 10.96 1.08 11.36 1.48 ;
      RECT 11.12 1.08 11.36 1.85 ;
      RECT 11.18 2.15 11.8 2.55 ;
      RECT 11.18 1.66 11.43 3.5 ;
      RECT 11.11 3.34 11.36 4.68 ;
      RECT 10.96 4.28 11.36 4.68 ;
  END
END UCL_DFF_LP

MACRO UCL_DFF_LP2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_LP2 0 0 ;
  SIZE 14.4 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 14.4 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.5 0.44 0.9 1.48 ;
        RECT 2.85 0.44 3.25 1.08 ;
        RECT 2.86 1.08 3.26 1.48 ;
        RECT 5.78 0.44 6.18 1.48 ;
        RECT 9.06 0.44 9.46 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 0 0.44 14.4 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 14.4 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.22 4.28 1.62 5.32 ;
        RECT 3.58 4.28 3.98 5.32 ;
        RECT 5.78 3.84 6.18 5.32 ;
        RECT 8.4 4.28 8.8 5.32 ;
        RECT 11.68 4.28 12.08 5.32 ;
        RECT 13.12 4.06 13.52 5.32 ;
        RECT 0 4.92 14.4 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 7.42 2.02 7.7 2.3 ;
      LAYER ME2 ;
        RECT 7.34 1.94 7.78 2.38 ;
      LAYER ME1 ;
        RECT 7.34 1.94 7.78 2.38 ;
        RECT 7.07 1.66 7.64 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9322 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025199 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME2 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME1 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.49 2.8 1.89 3.2 ;
        RECT 1.49 2.34 1.73 3.2 ;
        RECT 1.25 2.22 1.61 2.44 ;
        RECT 1.13 2.1 1.49 2.32 ;
        RECT 1.37 2.34 1.73 2.56 ;
        RECT 0.14 1.98 1.37 2.14 ;
        RECT 0.14 1.86 1.25 2.14 ;
        RECT 0.14 1.74 1.13 2.14 ;
        RECT 1.07 2.1 1.49 2.2 ;
        RECT 0.14 1.74 0.73 2.38 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 12.46 2.02 12.74 2.3 ;
      LAYER ME2 ;
        RECT 12.38 1.94 12.82 2.38 ;
      LAYER ME1 ;
        RECT 12.38 1.94 12.82 2.38 ;
        RECT 12.4 4.28 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.51 1.08 12.75 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1152 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 13.9 2.74 14.18 3.02 ;
      LAYER ME2 ;
        RECT 13.82 2.66 14.26 3.1 ;
      LAYER ME1 ;
        RECT 13.82 2.66 14.26 3.1 ;
        RECT 13.84 4.06 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 1.68 1.08 2.08 1.48 ;
      RECT 1.84 1.08 2.08 1.84 ;
      RECT 1.96 1.74 3.75 1.96 ;
      RECT 2.08 1.74 3.75 1.98 ;
      RECT 2.08 1.62 2.18 2.06 ;
      RECT 3.35 1.74 3.75 2.14 ;
      RECT 2.18 2.72 2.54 2.85 ;
      RECT 2.18 1.72 2.2 2.85 ;
      RECT 2.2 1.74 2.42 2.97 ;
      RECT 2.32 2.84 2.64 3.05 ;
      RECT 2.4 2.84 2.64 4.68 ;
      RECT 2.4 4.28 2.8 4.68 ;
      RECT 3.58 1.08 3.98 1.48 ;
      RECT 3.58 1.31 4.51 1.48 ;
      RECT 3.58 1.24 4.39 1.48 ;
      RECT 4.2 1.43 4.63 1.6 ;
      RECT 4.32 1.43 4.63 1.67 ;
      RECT 4.39 1.87 4.87 2.27 ;
      RECT 2.67 2.22 3.07 2.62 ;
      RECT 2.67 2.38 4.63 2.62 ;
      RECT 4.39 1.43 4.63 4.68 ;
      RECT 4.3 4.28 4.7 4.68 ;
      RECT 5.59 2.83 6 3.2 ;
      RECT 5.59 3.04 6.62 3.2 ;
      RECT 5.59 2.96 6.5 3.2 ;
      RECT 6.32 3.16 6.74 3.3 ;
      RECT 6.42 3.28 6.86 3.38 ;
      RECT 6.5 3.28 6.86 4.68 ;
      RECT 6.5 3.4 6.9 4.68 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.46 1.68 6.74 1.84 ;
      RECT 6.5 1.08 6.74 1.84 ;
      RECT 5.59 1.72 6.69 1.96 ;
      RECT 5.59 1.72 5.99 2.11 ;
      RECT 5.06 1.08 5.46 1.48 ;
      RECT 5.11 2.35 7.09 2.59 ;
      RECT 6.69 2.35 7.09 2.87 ;
      RECT 6.69 2.63 9.76 2.87 ;
      RECT 4.87 2.6 5.35 3 ;
      RECT 9.36 2.63 9.76 3.09 ;
      RECT 5.11 1.08 5.35 4.68 ;
      RECT 5.06 3.84 5.46 4.68 ;
      RECT 7.88 1.08 8.28 1.48 ;
      RECT 10.24 1.08 10.64 1.48 ;
      RECT 8.11 1.08 8.28 1.6 ;
      RECT 8.23 1.54 8.59 1.65 ;
      RECT 8.28 1.61 8.7 1.77 ;
      RECT 9.69 1.59 10.24 1.96 ;
      RECT 9.57 1.6 10.24 1.96 ;
      RECT 8.28 1.3 8.4 1.77 ;
      RECT 8.4 1.42 8.52 1.89 ;
      RECT 9.7 1.24 10.24 1.96 ;
      RECT 8.52 1.72 10.24 1.96 ;
      RECT 10 2.15 10.94 2.55 ;
      RECT 9.05 3.13 9.17 3.8 ;
      RECT 7.74 3.11 9.05 3.35 ;
      RECT 7.62 3.21 7.74 3.67 ;
      RECT 7.51 3.33 7.94 3.45 ;
      RECT 8.93 3.25 9.29 3.45 ;
      RECT 9.03 3.25 9.29 3.47 ;
      RECT 7.39 3.44 7.84 3.55 ;
      RECT 7.39 3.44 7.74 3.67 ;
      RECT 9.05 3.25 9.29 3.8 ;
      RECT 10 1.24 10.24 3.8 ;
      RECT 9.05 3.56 10.24 3.8 ;
      RECT 7.22 3.56 7.62 4.68 ;
      RECT 9.58 3.56 9.98 4.68 ;
      RECT 10.96 1.08 11.36 1.48 ;
      RECT 11.12 1.08 11.36 1.85 ;
      RECT 11.18 2.15 11.8 2.55 ;
      RECT 11.18 1.66 11.43 3.5 ;
      RECT 11.11 3.34 11.36 4.68 ;
      RECT 10.96 4.28 11.36 4.68 ;
  END
END UCL_DFF_LP2

MACRO UCL_DFF_LP4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_LP4 0 0 ;
  SIZE 15.12 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 15.12 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.5 0.44 0.9 1.48 ;
        RECT 2.85 0.44 3.25 1.08 ;
        RECT 2.86 1.08 3.26 1.48 ;
        RECT 5.78 0.44 6.18 1.48 ;
        RECT 9.06 0.44 9.46 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 0 0.44 15.12 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 15.12 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.22 4.28 1.62 5.32 ;
        RECT 3.58 4.28 3.98 5.32 ;
        RECT 5.78 3.84 6.18 5.32 ;
        RECT 8.4 4.28 8.8 5.32 ;
        RECT 11.68 4.28 12.08 5.32 ;
        RECT 13.12 4.06 13.52 5.32 ;
        RECT 14.56 4.06 14.96 5.32 ;
        RECT 0 4.92 15.12 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 7.42 2.02 7.7 2.3 ;
      LAYER ME2 ;
        RECT 7.34 1.94 7.78 2.38 ;
      LAYER ME1 ;
        RECT 7.34 1.94 7.78 2.38 ;
        RECT 7.07 1.66 7.64 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9322 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.025199 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME2 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME1 ;
      ANTENNAMAXAREACAR 5.885101 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 19.098478 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.49 2.8 1.89 3.2 ;
        RECT 1.49 2.34 1.73 3.2 ;
        RECT 1.25 2.22 1.61 2.44 ;
        RECT 1.13 2.1 1.49 2.32 ;
        RECT 1.37 2.34 1.73 2.56 ;
        RECT 0.14 1.98 1.37 2.14 ;
        RECT 0.14 1.86 1.25 2.14 ;
        RECT 0.14 1.74 1.13 2.14 ;
        RECT 1.07 2.1 1.49 2.2 ;
        RECT 0.14 1.74 0.73 2.38 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 12.46 2.02 12.74 2.3 ;
      LAYER ME2 ;
        RECT 12.38 1.94 12.82 2.38 ;
      LAYER ME1 ;
        RECT 12.38 1.94 12.82 2.38 ;
        RECT 12.4 4.28 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.51 1.08 12.75 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1152 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.7128 LAYER ME1 ;
    ANTENNADIFFAREA 0.7128 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 13.9 2.74 14.18 3.02 ;
      LAYER ME2 ;
        RECT 13.82 2.66 14.26 3.1 ;
      LAYER ME1 ;
        RECT 13.82 2.66 14.26 3.1 ;
        RECT 13.84 4.06 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
    END
  END Q
  OBS
    LAYER ME1 ;
      RECT 1.68 1.08 2.08 1.48 ;
      RECT 1.84 1.08 2.08 1.84 ;
      RECT 1.96 1.74 3.75 1.96 ;
      RECT 2.08 1.74 3.75 1.98 ;
      RECT 2.08 1.62 2.18 2.06 ;
      RECT 3.35 1.74 3.75 2.14 ;
      RECT 2.18 2.72 2.54 2.85 ;
      RECT 2.18 1.72 2.2 2.85 ;
      RECT 2.2 1.74 2.42 2.97 ;
      RECT 2.32 2.84 2.64 3.05 ;
      RECT 2.4 2.84 2.64 4.68 ;
      RECT 2.4 4.28 2.8 4.68 ;
      RECT 3.58 1.08 3.98 1.48 ;
      RECT 3.58 1.31 4.51 1.48 ;
      RECT 3.58 1.24 4.39 1.48 ;
      RECT 4.2 1.43 4.63 1.6 ;
      RECT 4.32 1.43 4.63 1.67 ;
      RECT 4.39 1.87 4.87 2.27 ;
      RECT 2.67 2.22 3.07 2.62 ;
      RECT 2.67 2.38 4.63 2.62 ;
      RECT 4.39 1.43 4.63 4.68 ;
      RECT 4.3 4.28 4.7 4.68 ;
      RECT 5.59 2.83 6 3.2 ;
      RECT 5.59 3.04 6.62 3.2 ;
      RECT 5.59 2.96 6.5 3.2 ;
      RECT 6.32 3.16 6.74 3.3 ;
      RECT 6.42 3.28 6.86 3.38 ;
      RECT 6.5 3.28 6.86 4.68 ;
      RECT 6.5 3.4 6.9 4.68 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.46 1.68 6.74 1.84 ;
      RECT 6.5 1.08 6.74 1.84 ;
      RECT 5.59 1.72 6.69 1.96 ;
      RECT 5.59 1.72 5.99 2.11 ;
      RECT 5.06 1.08 5.46 1.48 ;
      RECT 5.11 2.35 7.09 2.59 ;
      RECT 6.69 2.35 7.09 2.87 ;
      RECT 6.69 2.63 9.76 2.87 ;
      RECT 4.87 2.6 5.35 3 ;
      RECT 9.36 2.63 9.76 3.09 ;
      RECT 5.11 1.08 5.35 4.68 ;
      RECT 5.06 3.84 5.46 4.68 ;
      RECT 7.88 1.08 8.28 1.48 ;
      RECT 10.24 1.08 10.64 1.48 ;
      RECT 8.11 1.08 8.28 1.6 ;
      RECT 8.23 1.54 8.59 1.65 ;
      RECT 8.28 1.61 8.7 1.77 ;
      RECT 9.69 1.59 10.24 1.96 ;
      RECT 9.57 1.6 10.24 1.96 ;
      RECT 8.28 1.3 8.4 1.77 ;
      RECT 8.4 1.42 8.52 1.89 ;
      RECT 9.7 1.24 10.24 1.96 ;
      RECT 8.52 1.72 10.24 1.96 ;
      RECT 10 2.15 10.94 2.55 ;
      RECT 9.05 3.13 9.17 3.8 ;
      RECT 7.74 3.11 9.05 3.35 ;
      RECT 7.62 3.21 7.74 3.67 ;
      RECT 7.51 3.33 7.94 3.45 ;
      RECT 8.93 3.25 9.29 3.45 ;
      RECT 9.03 3.25 9.29 3.47 ;
      RECT 7.39 3.44 7.84 3.55 ;
      RECT 7.39 3.44 7.74 3.67 ;
      RECT 9.05 3.25 9.29 3.8 ;
      RECT 10 1.24 10.24 3.8 ;
      RECT 9.05 3.56 10.24 3.8 ;
      RECT 7.22 3.56 7.62 4.68 ;
      RECT 9.58 3.56 9.98 4.68 ;
      RECT 10.96 1.08 11.36 1.48 ;
      RECT 11.12 1.08 11.36 1.85 ;
      RECT 11.18 2.15 11.8 2.55 ;
      RECT 11.18 1.66 11.43 3.5 ;
      RECT 11.11 3.34 11.36 4.68 ;
      RECT 10.96 4.28 11.36 4.68 ;
  END
END UCL_DFF_LP4

MACRO UCL_DFF_RES
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_RES 0 0 ;
  SIZE 17.28 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 17.28 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.52 0.44 2.92 1.48 ;
        RECT 3.24 0.44 3.64 1.48 ;
        RECT 4.68 0.44 5.08 1.48 ;
        RECT 7.22 0.44 7.62 1.48 ;
        RECT 10.5 0.44 10.9 1.48 ;
        RECT 12.4 0.44 12.8 1.48 ;
        RECT 13.84 0.44 14.24 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 0 0.44 17.28 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 17.28 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 3.24 3.56 3.64 5.32 ;
        RECT 5.14 3.56 5.54 5.32 ;
        RECT 7.22 3.56 7.62 5.32 ;
        RECT 9.84 3.58 10.24 5.32 ;
        RECT 13.84 3.56 14.24 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 0 4.92 17.28 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 8.86 2.02 9.14 2.3 ;
      LAYER ME2 ;
        RECT 8.78 1.94 9.22 2.38 ;
      LAYER ME1 ;
        RECT 8.78 1.94 9.22 2.38 ;
        RECT 8.51 1.66 9.08 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.825 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.535882 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 2.518315 LAYER ME1 ;
      ANTENNAMAXAREACAR 2.518315 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 7.740786 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 7.740786 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.15 2.8 1.55 3.2 ;
        RECT 1.15 2.34 1.39 3.2 ;
        RECT 0.14 2.22 1.27 2.38 ;
        RECT 0.14 2.16 1.15 2.38 ;
        RECT 1.09 2.34 1.39 2.56 ;
        RECT 0.14 2.04 1.09 2.38 ;
        RECT 0.97 2.34 1.39 2.5 ;
        RECT 0.14 1.98 0.97 2.38 ;
        RECT 0.14 1.86 0.91 2.38 ;
        RECT 0.14 1.74 0.79 2.38 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 15.34 2.02 15.62 2.3 ;
      LAYER ME2 ;
        RECT 15.26 1.94 15.7 2.38 ;
      LAYER ME1 ;
        RECT 15.26 1.94 15.7 2.38 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.39 1.08 15.63 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 16.78 2.74 17.06 3.02 ;
      LAYER ME2 ;
        RECT 16.7 2.66 17.14 3.1 ;
      LAYER ME1 ;
        RECT 16.7 2.66 17.14 3.1 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.8 1.08 17.04 4.68 ;
    END
  END Q
  PIN RES
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.6984 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 4.97 2.74 5.25 3.02 ;
        RECT 13.64 2.74 13.92 3.02 ;
      LAYER ME2 ;
        RECT 4.89 2.84 14 3.12 ;
        RECT 13.56 2.66 14 3.12 ;
        RECT 4.89 2.66 5.62 3.12 ;
      LAYER ME1 ;
        RECT 13.56 2.66 14 3.1 ;
        RECT 4.89 2.66 5.33 3.1 ;
    END
  END RES
  OBS
    LAYER ME1 ;
      RECT 1.34 1.08 1.74 1.48 ;
      RECT 1.5 1.62 1.76 1.84 ;
      RECT 1.74 1.64 1.84 1.98 ;
      RECT 1.5 1.08 1.74 1.84 ;
      RECT 1.62 1.74 3.87 1.96 ;
      RECT 1.74 1.74 3.87 1.98 ;
      RECT 3.47 1.74 3.87 2.14 ;
      RECT 1.84 2.72 2.2 2.84 ;
      RECT 1.84 1.72 1.86 2.84 ;
      RECT 1.86 1.74 2.08 2.96 ;
      RECT 1.98 2.84 2.3 3.04 ;
      RECT 2.06 2.84 2.3 4.68 ;
      RECT 2.06 3.56 2.46 4.68 ;
      RECT 3.96 1.08 4.36 1.48 ;
      RECT 5.77 1.82 6.31 2.22 ;
      RECT 2.33 2.22 2.73 2.62 ;
      RECT 4.12 2.17 6.07 2.42 ;
      RECT 2.33 2.38 4.36 2.62 ;
      RECT 4.12 1.08 4.36 4.68 ;
      RECT 3.96 3.56 4.36 4.68 ;
      RECT 7.03 2.83 7.43 3.2 ;
      RECT 7.03 3.04 8.06 3.2 ;
      RECT 7.03 2.96 7.94 3.2 ;
      RECT 7.76 3.16 8.18 3.3 ;
      RECT 7.86 3.16 8.18 3.38 ;
      RECT 7.94 3.16 8.18 4.68 ;
      RECT 7.94 3.56 8.34 4.68 ;
      RECT 7.94 1.08 8.34 1.48 ;
      RECT 7.91 1.69 8.18 1.84 ;
      RECT 7.94 1.08 8.18 1.84 ;
      RECT 7.03 1.72 8.13 1.96 ;
      RECT 7.03 1.72 7.43 2.11 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.55 2.35 8.53 2.59 ;
      RECT 8.13 2.35 8.53 2.86 ;
      RECT 8.13 2.62 11.2 2.86 ;
      RECT 10.6 2.62 11.2 2.98 ;
      RECT 6.31 2.6 6.79 3 ;
      RECT 10.72 2.62 11.2 3.06 ;
      RECT 10.8 2.62 11.2 3.09 ;
      RECT 6.55 1.08 6.79 4.68 ;
      RECT 6.5 3.56 6.9 4.68 ;
      RECT 9.32 1.08 9.72 1.48 ;
      RECT 11.68 1.08 12.08 1.48 ;
      RECT 9.56 1.08 9.72 1.6 ;
      RECT 9.68 1.54 10.04 1.64 ;
      RECT 9.72 1.62 10.14 1.76 ;
      RECT 11.01 1.6 11.68 1.96 ;
      RECT 9.72 1.3 9.84 1.76 ;
      RECT 11.13 1.58 11.68 1.96 ;
      RECT 9.84 1.72 11.68 1.88 ;
      RECT 9.84 1.42 9.96 1.88 ;
      RECT 11.15 1.24 11.68 1.96 ;
      RECT 9.96 1.82 12.85 1.96 ;
      RECT 11.44 1.82 12.85 2.06 ;
      RECT 12.45 1.74 12.85 2.14 ;
      RECT 9.3 3.1 10.58 3.34 ;
      RECT 9.06 3.27 9.45 3.44 ;
      RECT 9.18 3.15 9.3 3.61 ;
      RECT 9.01 3.39 9.45 3.44 ;
      RECT 10.36 3.34 10.82 3.44 ;
      RECT 10.46 3.34 10.82 3.56 ;
      RECT 8.89 3.44 9.35 3.49 ;
      RECT 8.89 3.44 9.3 3.61 ;
      RECT 10.46 3.46 10.92 3.56 ;
      RECT 11.44 1.24 11.68 3.8 ;
      RECT 10.58 3.22 10.7 3.68 ;
      RECT 8.66 3.56 9.18 3.73 ;
      RECT 10.7 3.56 11.68 3.8 ;
      RECT 8.66 3.56 9.06 4.68 ;
      RECT 11.02 3.56 11.42 4.68 ;
      RECT 13.12 1.08 13.52 1.48 ;
      RECT 12.98 2.27 14.68 2.39 ;
      RECT 13.2 2.15 14.68 2.39 ;
      RECT 13.2 1.08 13.44 2.44 ;
      RECT 13.1 2.17 13.2 2.73 ;
      RECT 12.86 2.39 13.39 2.51 ;
      RECT 14.28 2.15 14.68 2.55 ;
      RECT 12.74 2.51 13.32 2.63 ;
      RECT 12.74 2.51 13.1 2.85 ;
      RECT 12.74 2.51 12.98 4.68 ;
      RECT 12.66 3.56 13.06 4.68 ;
  END
END UCL_DFF_RES

MACRO UCL_DFF_RES2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_RES2 0 0 ;
  SIZE 18 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 8.51 1.66 9.08 2.07 ;
        RECT 8.78 1.94 9.22 2.38 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.74 0.79 2.38 ;
        RECT 0.14 1.86 0.91 2.38 ;
        RECT 0.14 1.98 0.97 2.38 ;
        RECT 0.97 2.34 1.39 2.5 ;
        RECT 0.14 2.04 1.09 2.38 ;
        RECT 1.09 2.34 1.39 2.56 ;
        RECT 0.14 2.16 1.15 2.38 ;
        RECT 0.14 2.22 1.27 2.38 ;
        RECT 1.15 2.34 1.39 3.2 ;
        RECT 1.15 2.8 1.55 3.2 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 15.39 1.08 15.63 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.28 3.56 15.68 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 16.8 1.08 17.04 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.72 3.56 17.12 4.68 ;
    END
  END Q
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 18 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.52 0.44 2.92 1.48 ;
        RECT 3.24 0.44 3.64 1.48 ;
        RECT 4.68 0.44 5.08 1.48 ;
        RECT 7.22 0.44 7.62 1.48 ;
        RECT 10.5 0.44 10.9 1.48 ;
        RECT 12.4 0.44 12.8 1.48 ;
        RECT 13.84 0.44 14.24 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 0 0.44 18 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 18 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 3.24 3.56 3.64 5.32 ;
        RECT 5.14 3.56 5.54 5.32 ;
        RECT 7.22 3.56 7.62 5.32 ;
        RECT 9.84 3.58 10.24 5.32 ;
        RECT 13.84 3.56 14.24 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 0 4.92 18 5.32 ;
    END
  END vddd
  PIN RES
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.6984 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 4.97 2.74 5.25 3.02 ;
        RECT 13.64 2.74 13.92 3.02 ;
      LAYER ME1 ;
        RECT 13.56 2.66 14 3.1 ;
        RECT 4.89 2.66 5.33 3.1 ;
      LAYER ME2 ;
        RECT 4.89 2.84 14 3.12 ;
        RECT 13.56 2.66 14 3.12 ;
        RECT 4.89 2.66 5.62 3.12 ;
    END
  END RES
  OBS
    LAYER ME1 ;
      RECT 1.34 1.08 1.74 1.48 ;
      RECT 1.5 1.62 1.76 1.84 ;
      RECT 1.74 1.64 1.84 1.98 ;
      RECT 1.5 1.08 1.74 1.84 ;
      RECT 1.62 1.74 3.87 1.96 ;
      RECT 1.74 1.74 3.87 1.98 ;
      RECT 3.47 1.74 3.87 2.14 ;
      RECT 1.84 2.72 2.2 2.84 ;
      RECT 1.84 1.72 1.86 2.84 ;
      RECT 1.86 1.74 2.08 2.96 ;
      RECT 1.98 2.84 2.3 3.04 ;
      RECT 2.06 2.84 2.3 4.68 ;
      RECT 2.06 3.56 2.46 4.68 ;
      RECT 3.96 1.08 4.36 1.48 ;
      RECT 5.77 1.82 6.31 2.22 ;
      RECT 2.33 2.22 2.73 2.62 ;
      RECT 4.12 2.17 6.07 2.42 ;
      RECT 2.33 2.38 4.36 2.62 ;
      RECT 4.12 1.08 4.36 4.68 ;
      RECT 3.96 3.56 4.36 4.68 ;
      RECT 7.03 2.83 7.43 3.2 ;
      RECT 7.03 3.04 8.06 3.2 ;
      RECT 7.03 2.96 7.94 3.2 ;
      RECT 7.76 3.16 8.18 3.3 ;
      RECT 7.86 3.16 8.18 3.38 ;
      RECT 7.94 3.16 8.18 4.68 ;
      RECT 7.94 3.56 8.34 4.68 ;
      RECT 7.94 1.08 8.34 1.48 ;
      RECT 7.91 1.69 8.18 1.84 ;
      RECT 7.94 1.08 8.18 1.84 ;
      RECT 7.03 1.72 8.13 1.96 ;
      RECT 7.03 1.72 7.43 2.11 ;
      RECT 6.5 1.08 6.9 1.48 ;
      RECT 6.55 2.35 8.53 2.59 ;
      RECT 8.13 2.35 8.53 2.86 ;
      RECT 8.13 2.62 11.2 2.86 ;
      RECT 10.6 2.62 11.2 2.98 ;
      RECT 6.31 2.6 6.79 3 ;
      RECT 10.72 2.62 11.2 3.06 ;
      RECT 10.8 2.62 11.2 3.09 ;
      RECT 6.55 1.08 6.79 4.68 ;
      RECT 6.5 3.56 6.9 4.68 ;
      RECT 9.32 1.08 9.72 1.48 ;
      RECT 11.68 1.08 12.08 1.48 ;
      RECT 9.56 1.08 9.72 1.6 ;
      RECT 9.68 1.54 10.04 1.64 ;
      RECT 9.72 1.62 10.14 1.76 ;
      RECT 11.01 1.6 11.68 1.96 ;
      RECT 9.72 1.3 9.84 1.76 ;
      RECT 11.13 1.58 11.68 1.96 ;
      RECT 9.84 1.72 11.68 1.88 ;
      RECT 9.84 1.42 9.96 1.88 ;
      RECT 11.15 1.24 11.68 1.96 ;
      RECT 9.96 1.82 12.85 1.96 ;
      RECT 11.44 1.82 12.85 2.06 ;
      RECT 12.45 1.74 12.85 2.14 ;
      RECT 9.3 3.1 10.58 3.34 ;
      RECT 9.06 3.27 9.45 3.44 ;
      RECT 9.18 3.15 9.3 3.61 ;
      RECT 9.01 3.39 9.45 3.44 ;
      RECT 10.36 3.34 10.82 3.44 ;
      RECT 10.46 3.34 10.82 3.56 ;
      RECT 8.89 3.44 9.35 3.49 ;
      RECT 8.89 3.44 9.3 3.61 ;
      RECT 10.46 3.46 10.92 3.56 ;
      RECT 11.44 1.24 11.68 3.8 ;
      RECT 10.58 3.22 10.7 3.68 ;
      RECT 8.66 3.56 9.18 3.73 ;
      RECT 10.7 3.56 11.68 3.8 ;
      RECT 8.66 3.56 9.06 4.68 ;
      RECT 11.02 3.56 11.42 4.68 ;
      RECT 13.12 1.08 13.52 1.48 ;
      RECT 12.98 2.27 14.68 2.39 ;
      RECT 13.2 2.15 14.68 2.39 ;
      RECT 13.2 1.08 13.44 2.44 ;
      RECT 13.1 2.17 13.2 2.73 ;
      RECT 12.86 2.39 13.39 2.51 ;
      RECT 14.28 2.15 14.68 2.55 ;
      RECT 12.74 2.51 13.32 2.63 ;
      RECT 12.74 2.51 13.1 2.85 ;
      RECT 12.74 2.51 12.98 4.68 ;
      RECT 12.66 3.56 13.06 4.68 ;
  END
END UCL_DFF_RES2

MACRO UCL_DFF_SCAN
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_SCAN 0 0 ;
  SIZE 18.72 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.16 4.28 18.56 4.68 ;
        RECT 18.14 2.66 18.58 3.1 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 16.83 1.08 17.07 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.72 4.28 17.12 4.68 ;
        RECT 16.7 1.94 17.14 2.38 ;
    END
  END Q
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 18.72 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.4 0.44 1.8 1.48 ;
        RECT 3.76 0.44 4.16 1.48 ;
        RECT 4.82 0.44 5.22 1.48 ;
        RECT 7.17 0.44 7.57 1.08 ;
        RECT 7.18 1.08 7.58 1.48 ;
        RECT 10.1 0.44 10.5 1.48 ;
        RECT 13.38 0.44 13.78 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 0 0.44 18.72 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 18.72 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.4 3.56 1.8 5.32 ;
        RECT 3.76 3.56 4.16 5.32 ;
        RECT 5.54 4.28 5.94 5.32 ;
        RECT 7.9 4.28 8.3 5.32 ;
        RECT 10.1 3.84 10.5 5.32 ;
        RECT 12.72 4.28 13.12 5.32 ;
        RECT 16 4.28 16.4 5.32 ;
        RECT 17.44 4.28 17.84 5.32 ;
        RECT 0 4.92 18.72 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.634259 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.777778 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 11.74 2.02 12.02 2.3 ;
      LAYER ME1 ;
        RECT 11.66 1.94 12.1 2.38 ;
        RECT 11.39 1.66 11.96 2.07 ;
      LAYER ME2 ;
        RECT 11.66 1.94 12.1 2.38 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3124 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.104 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.02 1.94 2.3 ;
      LAYER ME1 ;
        RECT 1.58 1.94 2.29 2.38 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.02 2.38 ;
    END
  END D
  PIN SCAN_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1484 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.928 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME1 ;
        RECT 0.14 2.66 2.75 3.1 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END SCAN_EN
  PIN SCAN_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0464 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.82 2.74 4.1 3.02 ;
      LAYER ME1 ;
        RECT 3.53 2.66 4.18 3.1 ;
      LAYER ME2 ;
        RECT 3.74 2.66 4.18 3.1 ;
    END
  END SCAN_IN
  OBS
    LAYER ME1 ;
      RECT 0.14 3.56 1.08 4.46 ;
      RECT 0.68 3.56 1.08 4.68 ;
      RECT 0.14 1.08 1.08 1.48 ;
      RECT 2.58 1.08 2.98 1.48 ;
      RECT 2.74 1.08 2.98 2.07 ;
      RECT 3.92 1.9 5.57 2.14 ;
      RECT 5.05 1.74 5.45 2.14 ;
      RECT 2.86 1.94 4.16 2.18 ;
      RECT 2.86 1.94 3.46 2.19 ;
      RECT 2.98 1.85 2.99 2.2 ;
      RECT 5.39 2.1 5.81 2.2 ;
      RECT 5.45 1.86 5.57 2.32 ;
      RECT 5.57 2.22 5.93 2.44 ;
      RECT 2.99 1.94 3.46 2.38 ;
      RECT 5.57 1.98 5.69 2.44 ;
      RECT 5.69 2.1 5.81 2.56 ;
      RECT 5.81 2.34 6.05 3.2 ;
      RECT 5.81 2.8 6.21 3.2 ;
      RECT 2.99 1.94 3.23 3.38 ;
      RECT 2.91 3.25 2.98 4.68 ;
      RECT 2.79 3.32 3.19 3.5 ;
      RECT 2.98 3.24 2.99 3.59 ;
      RECT 2.67 3.44 3.07 3.58 ;
      RECT 2.99 1.86 3.07 3.58 ;
      RECT 2.58 3.56 2.98 4.68 ;
      RECT 6 1.08 6.4 1.48 ;
      RECT 6.16 1.08 6.4 1.84 ;
      RECT 6.28 1.74 8.07 1.96 ;
      RECT 6.4 1.74 8.07 1.98 ;
      RECT 6.4 1.62 6.5 2.06 ;
      RECT 7.67 1.74 8.07 2.14 ;
      RECT 6.5 2.72 6.86 2.85 ;
      RECT 6.5 1.72 6.52 2.85 ;
      RECT 6.52 1.74 6.74 2.97 ;
      RECT 6.64 2.84 6.96 3.05 ;
      RECT 6.72 2.84 6.96 4.68 ;
      RECT 6.72 4.28 7.12 4.68 ;
      RECT 7.9 1.08 8.3 1.48 ;
      RECT 7.9 1.31 8.83 1.48 ;
      RECT 7.9 1.24 8.71 1.48 ;
      RECT 8.52 1.43 8.95 1.6 ;
      RECT 8.64 1.43 8.95 1.67 ;
      RECT 8.71 1.87 9.19 2.27 ;
      RECT 6.99 2.22 7.39 2.62 ;
      RECT 6.99 2.38 8.95 2.62 ;
      RECT 8.71 1.43 8.95 4.68 ;
      RECT 8.62 4.28 9.02 4.68 ;
      RECT 9.91 2.83 10.32 3.2 ;
      RECT 9.91 3.04 10.94 3.2 ;
      RECT 9.91 2.96 10.82 3.2 ;
      RECT 10.64 3.16 11.06 3.3 ;
      RECT 10.74 3.28 11.18 3.38 ;
      RECT 10.82 3.28 11.18 4.68 ;
      RECT 10.82 3.4 11.22 4.68 ;
      RECT 10.82 1.08 11.22 1.48 ;
      RECT 10.78 1.68 11.06 1.84 ;
      RECT 10.82 1.08 11.06 1.84 ;
      RECT 9.91 1.72 11.01 1.96 ;
      RECT 9.91 1.72 10.31 2.11 ;
      RECT 9.38 1.08 9.78 1.48 ;
      RECT 9.43 2.35 11.41 2.59 ;
      RECT 11.01 2.35 11.41 2.87 ;
      RECT 11.01 2.63 14.08 2.87 ;
      RECT 9.19 2.6 9.67 3 ;
      RECT 13.68 2.63 14.08 3.09 ;
      RECT 9.43 1.08 9.67 4.68 ;
      RECT 9.38 3.84 9.78 4.68 ;
      RECT 12.2 1.08 12.6 1.48 ;
      RECT 14.56 1.08 14.96 1.48 ;
      RECT 12.43 1.08 12.6 1.6 ;
      RECT 12.55 1.54 12.91 1.65 ;
      RECT 12.6 1.61 13.02 1.77 ;
      RECT 14.01 1.59 14.56 1.96 ;
      RECT 13.89 1.6 14.56 1.96 ;
      RECT 12.6 1.3 12.72 1.77 ;
      RECT 12.72 1.42 12.84 1.89 ;
      RECT 14.02 1.24 14.56 1.96 ;
      RECT 12.84 1.72 14.56 1.96 ;
      RECT 14.32 2.15 15.26 2.55 ;
      RECT 13.37 3.13 13.49 3.8 ;
      RECT 12.06 3.11 13.37 3.35 ;
      RECT 11.94 3.21 12.06 3.67 ;
      RECT 11.83 3.33 12.26 3.45 ;
      RECT 13.25 3.25 13.61 3.45 ;
      RECT 13.35 3.25 13.61 3.47 ;
      RECT 11.71 3.44 12.16 3.55 ;
      RECT 11.71 3.44 12.06 3.67 ;
      RECT 13.37 3.25 13.61 3.8 ;
      RECT 14.32 1.24 14.56 3.8 ;
      RECT 13.37 3.56 14.56 3.8 ;
      RECT 11.54 3.56 11.94 4.68 ;
      RECT 13.9 3.56 14.3 4.68 ;
      RECT 15.28 1.08 15.68 1.48 ;
      RECT 15.44 1.08 15.68 1.85 ;
      RECT 15.5 2.15 16.12 2.55 ;
      RECT 15.5 1.66 15.75 3.5 ;
      RECT 15.43 3.34 15.68 4.68 ;
      RECT 15.28 4.28 15.68 4.68 ;
    LAYER ME2 ;
      RECT 3.02 1.94 3.46 2.38 ;
  END
END UCL_DFF_SCAN

MACRO UCL_DFF_SET
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_SET 0 0 ;
  SIZE 18.72 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 18.72 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.96 0.44 4.36 1.48 ;
        RECT 4.68 0.44 5.08 1.48 ;
        RECT 6.12 0.44 6.52 1.48 ;
        RECT 8.66 0.44 9.06 1.48 ;
        RECT 11.94 0.44 12.34 1.48 ;
        RECT 13.84 0.44 14.24 1.48 ;
        RECT 15.28 0.44 15.68 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 0 0.44 18.72 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 18.72 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 4.68 3.56 5.08 5.32 ;
        RECT 6.58 3.56 6.98 5.32 ;
        RECT 8.66 3.56 9.06 5.32 ;
        RECT 11.28 3.58 11.68 5.32 ;
        RECT 15.28 3.56 15.68 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 0 4.92 18.72 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.3883 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3728 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.185287 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.190476 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 10.3 2.02 10.58 2.3 ;
      LAYER ME2 ;
        RECT 10.22 1.94 10.66 2.38 ;
      LAYER ME1 ;
        RECT 10.22 1.94 10.66 2.38 ;
        RECT 9.95 1.66 10.52 2.07 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 18.22 2.74 18.5 3.02 ;
      LAYER ME2 ;
        RECT 18.14 2.66 18.58 3.1 ;
      LAYER ME1 ;
        RECT 18.14 2.66 18.58 3.1 ;
        RECT 18.16 3.56 18.56 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.24 1.08 18.48 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 16.78 2.02 17.06 2.3 ;
      LAYER ME2 ;
        RECT 16.7 1.94 17.14 2.38 ;
      LAYER ME1 ;
        RECT 16.7 1.94 17.14 2.38 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.83 1.08 17.07 4.68 ;
    END
  END Q
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.6984 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 6.41 2.74 6.69 3.02 ;
        RECT 15.08 2.74 15.36 3.02 ;
      LAYER ME2 ;
        RECT 6.33 2.84 15.44 3.12 ;
        RECT 15 2.66 15.44 3.12 ;
        RECT 6.33 2.66 7.06 3.12 ;
      LAYER ME1 ;
        RECT 15 2.66 15.44 3.1 ;
        RECT 6.33 2.66 6.77 3.1 ;
    END
  END SET
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.96 1.74 2.23 2.38 ;
      RECT 0.96 1.86 2.35 2.38 ;
      RECT 0.86 1.94 2.35 2.38 ;
      RECT 0.86 2.22 2.71 2.38 ;
      RECT 0.86 1.98 2.41 2.38 ;
      RECT 2.41 2.04 2.53 2.5 ;
      RECT 2.53 2.16 2.59 2.56 ;
      RECT 2.59 2.34 2.83 3.2 ;
      RECT 2.59 2.8 2.99 3.2 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.78 1.08 3.18 1.48 ;
      RECT 2.94 1.62 3.2 1.84 ;
      RECT 3.18 1.64 3.28 1.98 ;
      RECT 2.94 1.08 3.18 1.84 ;
      RECT 3.06 1.74 5.31 1.96 ;
      RECT 3.18 1.74 5.31 1.98 ;
      RECT 4.91 1.74 5.31 2.14 ;
      RECT 3.28 2.72 3.64 2.84 ;
      RECT 3.28 1.72 3.3 2.84 ;
      RECT 3.3 1.74 3.52 2.96 ;
      RECT 3.42 2.84 3.74 3.04 ;
      RECT 3.5 2.84 3.74 4.68 ;
      RECT 3.5 3.56 3.9 4.68 ;
      RECT 5.4 1.08 5.8 1.48 ;
      RECT 7.21 1.82 7.75 2.22 ;
      RECT 3.77 2.22 4.17 2.62 ;
      RECT 5.56 2.17 7.51 2.42 ;
      RECT 3.77 2.38 5.8 2.62 ;
      RECT 5.56 1.08 5.8 4.68 ;
      RECT 5.4 3.56 5.8 4.68 ;
      RECT 8.47 2.83 8.87 3.2 ;
      RECT 8.47 3.04 9.5 3.2 ;
      RECT 8.47 2.96 9.38 3.2 ;
      RECT 9.2 3.16 9.62 3.3 ;
      RECT 9.3 3.16 9.62 3.38 ;
      RECT 9.38 3.16 9.62 4.68 ;
      RECT 9.38 3.56 9.78 4.68 ;
      RECT 9.38 1.08 9.78 1.48 ;
      RECT 9.35 1.69 9.62 1.84 ;
      RECT 9.38 1.08 9.62 1.84 ;
      RECT 8.47 1.72 9.57 1.96 ;
      RECT 8.47 1.72 8.87 2.11 ;
      RECT 7.94 1.08 8.34 1.48 ;
      RECT 7.99 2.35 9.97 2.59 ;
      RECT 9.57 2.35 9.97 2.86 ;
      RECT 9.57 2.62 12.64 2.86 ;
      RECT 12.04 2.62 12.64 2.98 ;
      RECT 7.75 2.6 8.23 3 ;
      RECT 12.16 2.62 12.64 3.06 ;
      RECT 12.24 2.62 12.64 3.09 ;
      RECT 7.99 1.08 8.23 4.68 ;
      RECT 7.94 3.56 8.34 4.68 ;
      RECT 10.76 1.08 11.16 1.48 ;
      RECT 13.12 1.08 13.52 1.48 ;
      RECT 11 1.08 11.16 1.6 ;
      RECT 11.12 1.54 11.48 1.64 ;
      RECT 11.16 1.62 11.58 1.76 ;
      RECT 12.45 1.6 13.12 1.96 ;
      RECT 11.16 1.3 11.28 1.76 ;
      RECT 12.57 1.58 13.12 1.96 ;
      RECT 11.28 1.72 13.12 1.88 ;
      RECT 11.28 1.42 11.4 1.88 ;
      RECT 12.59 1.24 13.12 1.96 ;
      RECT 11.4 1.82 14.29 1.96 ;
      RECT 12.88 1.82 14.29 2.06 ;
      RECT 13.89 1.74 14.29 2.14 ;
      RECT 10.74 3.1 12.02 3.34 ;
      RECT 10.5 3.27 10.89 3.44 ;
      RECT 10.62 3.15 10.74 3.61 ;
      RECT 10.45 3.39 10.89 3.44 ;
      RECT 11.8 3.34 12.26 3.44 ;
      RECT 11.9 3.34 12.26 3.56 ;
      RECT 10.33 3.44 10.79 3.49 ;
      RECT 10.33 3.44 10.74 3.61 ;
      RECT 11.9 3.46 12.36 3.56 ;
      RECT 12.88 1.24 13.12 3.8 ;
      RECT 12.02 3.22 12.14 3.68 ;
      RECT 10.1 3.56 10.62 3.73 ;
      RECT 12.14 3.56 13.12 3.8 ;
      RECT 10.1 3.56 10.5 4.68 ;
      RECT 12.46 3.56 12.86 4.68 ;
      RECT 14.56 1.08 14.96 1.48 ;
      RECT 14.42 2.27 16.12 2.39 ;
      RECT 14.64 2.15 16.12 2.39 ;
      RECT 14.64 1.08 14.88 2.44 ;
      RECT 14.54 2.17 14.64 2.73 ;
      RECT 14.3 2.39 14.83 2.51 ;
      RECT 15.72 2.15 16.12 2.55 ;
      RECT 14.18 2.51 14.76 2.63 ;
      RECT 14.18 2.51 14.54 2.85 ;
      RECT 14.18 2.51 14.42 4.68 ;
      RECT 14.1 3.56 14.5 4.68 ;
  END
END UCL_DFF_SET

MACRO UCL_DFF_SET2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_DFF_SET2 0 0 ;
  SIZE 19.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 9.95 1.66 10.52 2.07 ;
        RECT 10.22 1.94 10.66 2.38 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END D
  PIN NQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.16 3.56 18.56 4.68 ;
    END
  END NQ
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 16.83 1.08 17.07 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.72 3.56 17.12 4.68 ;
    END
  END Q
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 18.72 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.96 0.44 4.36 1.48 ;
        RECT 4.68 0.44 5.08 1.48 ;
        RECT 6.12 0.44 6.52 1.48 ;
        RECT 8.66 0.44 9.06 1.48 ;
        RECT 11.94 0.44 12.34 1.48 ;
        RECT 13.84 0.44 14.24 1.48 ;
        RECT 15.28 0.44 15.68 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 0 0.44 18.72 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 18.72 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 4.68 3.56 5.08 5.32 ;
        RECT 6.58 3.56 6.98 5.32 ;
        RECT 8.66 3.56 9.06 5.32 ;
        RECT 11.28 3.58 11.68 5.32 ;
        RECT 15.28 3.56 15.68 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 0 4.92 18.72 5.32 ;
    END
  END vddd
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.6984 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 6.41 2.74 6.69 3.02 ;
        RECT 15.08 2.74 15.36 3.02 ;
      LAYER ME1 ;
        RECT 15 2.66 15.44 3.1 ;
        RECT 6.33 2.66 6.77 3.1 ;
      LAYER ME2 ;
        RECT 6.33 2.84 15.44 3.12 ;
        RECT 15 2.66 15.44 3.12 ;
        RECT 6.33 2.66 7.06 3.12 ;
    END
  END SET
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.96 1.74 2.23 2.38 ;
      RECT 0.96 1.86 2.35 2.38 ;
      RECT 0.86 1.94 2.35 2.38 ;
      RECT 0.86 2.22 2.71 2.38 ;
      RECT 0.86 1.98 2.41 2.38 ;
      RECT 2.41 2.04 2.53 2.5 ;
      RECT 2.53 2.16 2.59 2.56 ;
      RECT 2.59 2.34 2.83 3.2 ;
      RECT 2.59 2.8 2.99 3.2 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.78 1.08 3.18 1.48 ;
      RECT 2.94 1.62 3.2 1.84 ;
      RECT 3.18 1.64 3.28 1.98 ;
      RECT 2.94 1.08 3.18 1.84 ;
      RECT 3.06 1.74 5.31 1.96 ;
      RECT 3.18 1.74 5.31 1.98 ;
      RECT 4.91 1.74 5.31 2.14 ;
      RECT 3.28 2.72 3.64 2.84 ;
      RECT 3.28 1.72 3.3 2.84 ;
      RECT 3.3 1.74 3.52 2.96 ;
      RECT 3.42 2.84 3.74 3.04 ;
      RECT 3.5 2.84 3.74 4.68 ;
      RECT 3.5 3.56 3.9 4.68 ;
      RECT 5.4 1.08 5.8 1.48 ;
      RECT 7.21 1.82 7.75 2.22 ;
      RECT 3.77 2.22 4.17 2.62 ;
      RECT 5.56 2.17 7.51 2.42 ;
      RECT 3.77 2.38 5.8 2.62 ;
      RECT 5.56 1.08 5.8 4.68 ;
      RECT 5.4 3.56 5.8 4.68 ;
      RECT 8.47 2.83 8.87 3.2 ;
      RECT 8.47 3.04 9.5 3.2 ;
      RECT 8.47 2.96 9.38 3.2 ;
      RECT 9.2 3.16 9.62 3.3 ;
      RECT 9.3 3.16 9.62 3.38 ;
      RECT 9.38 3.16 9.62 4.68 ;
      RECT 9.38 3.56 9.78 4.68 ;
      RECT 9.38 1.08 9.78 1.48 ;
      RECT 9.35 1.69 9.62 1.84 ;
      RECT 9.38 1.08 9.62 1.84 ;
      RECT 8.47 1.72 9.57 1.96 ;
      RECT 8.47 1.72 8.87 2.11 ;
      RECT 7.94 1.08 8.34 1.48 ;
      RECT 7.99 2.35 9.97 2.59 ;
      RECT 9.57 2.35 9.97 2.86 ;
      RECT 9.57 2.62 12.64 2.86 ;
      RECT 12.04 2.62 12.64 2.98 ;
      RECT 7.75 2.6 8.23 3 ;
      RECT 12.16 2.62 12.64 3.06 ;
      RECT 12.24 2.62 12.64 3.09 ;
      RECT 7.99 1.08 8.23 4.68 ;
      RECT 7.94 3.56 8.34 4.68 ;
      RECT 10.76 1.08 11.16 1.48 ;
      RECT 13.12 1.08 13.52 1.48 ;
      RECT 11 1.08 11.16 1.6 ;
      RECT 11.12 1.54 11.48 1.64 ;
      RECT 11.16 1.62 11.58 1.76 ;
      RECT 12.45 1.6 13.12 1.96 ;
      RECT 11.16 1.3 11.28 1.76 ;
      RECT 12.57 1.58 13.12 1.96 ;
      RECT 11.28 1.72 13.12 1.88 ;
      RECT 11.28 1.42 11.4 1.88 ;
      RECT 12.59 1.24 13.12 1.96 ;
      RECT 11.4 1.82 14.29 1.96 ;
      RECT 12.88 1.82 14.29 2.06 ;
      RECT 13.89 1.74 14.29 2.14 ;
      RECT 10.74 3.1 12.02 3.34 ;
      RECT 10.5 3.27 10.89 3.44 ;
      RECT 10.62 3.15 10.74 3.61 ;
      RECT 10.45 3.39 10.89 3.44 ;
      RECT 11.8 3.34 12.26 3.44 ;
      RECT 11.9 3.34 12.26 3.56 ;
      RECT 10.33 3.44 10.79 3.49 ;
      RECT 10.33 3.44 10.74 3.61 ;
      RECT 11.9 3.46 12.36 3.56 ;
      RECT 12.88 1.24 13.12 3.8 ;
      RECT 12.02 3.22 12.14 3.68 ;
      RECT 10.1 3.56 10.62 3.73 ;
      RECT 12.14 3.56 13.12 3.8 ;
      RECT 10.1 3.56 10.5 4.68 ;
      RECT 12.46 3.56 12.86 4.68 ;
      RECT 14.56 1.08 14.96 1.48 ;
      RECT 14.42 2.27 16.45 2.39 ;
      RECT 14.64 2.15 16.45 2.39 ;
      RECT 14.64 1.08 14.88 2.44 ;
      RECT 14.54 2.17 14.64 2.73 ;
      RECT 14.3 2.39 14.83 2.51 ;
      RECT 16.05 2.15 16.45 2.55 ;
      RECT 14.18 2.51 14.76 2.63 ;
      RECT 14.18 2.51 14.54 2.85 ;
      RECT 14.18 2.51 14.42 4.68 ;
      RECT 14.1 3.56 14.5 4.68 ;
  END
END UCL_DFF_SET2

MACRO UCL_FA
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_FA 0 0 ;
  SIZE 11.52 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 11.52 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 3.76 0.44 4.16 1.48 ;
        RECT 5.2 0.44 5.6 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 0 0.44 11.52 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 11.52 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.84 1.28 5.32 ;
        RECT 3.76 3.84 4.16 5.32 ;
        RECT 5.2 3.84 5.6 5.32 ;
        RECT 6.64 3.84 7.04 5.32 ;
        RECT 10.24 4.06 10.64 5.32 ;
        RECT 0 4.92 11.52 5.32 ;
    END
  END vddd
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4852 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.76 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9504 LAYER ME1 ;
      ANTENNAGATEAREA 0.9504 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.56271 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.56271 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 6.060606 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 6.060606 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.082492 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.082492 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.12 3.32 3.4 3.6 ;
      LAYER ME2 ;
        RECT 3.04 3.24 3.48 3.68 ;
      LAYER ME1 ;
        RECT 2.81 3.36 5.67 3.6 ;
        RECT 5.27 3.34 5.67 3.6 ;
        RECT 3.04 3.24 3.48 3.68 ;
        RECT 2.08 3.2 3.21 3.44 ;
        RECT 2.08 2.88 2.32 3.44 ;
        RECT 0.65 2.88 2.32 3.12 ;
        RECT 0.65 2.72 1.05 3.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6808 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5952 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9504 LAYER ME1 ;
      ANTENNAGATEAREA 0.9504 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.768519 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.768519 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 6.939394 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 6.939394 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.082492 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.082492 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.68 1.83 3.96 2.11 ;
      LAYER ME2 ;
        RECT 3.6 1.75 4.04 2.19 ;
      LAYER ME1 ;
        RECT 6.86 1.72 7.26 2.04 ;
        RECT 5.05 1.75 7.26 1.99 ;
        RECT 3.11 1.91 5.29 2 ;
        RECT 3.53 1.76 7.26 1.99 ;
        RECT 3.6 1.75 4.04 2.19 ;
        RECT 3.53 1.75 4.04 2.15 ;
        RECT 3.11 1.91 4.04 2.15 ;
        RECT 2.09 2.04 3.35 2.28 ;
        RECT 1.37 2.2 2.33 2.44 ;
        RECT 1.37 2.2 1.77 2.6 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7096 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.88 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.7128 LAYER ME1 ;
      ANTENNAGATEAREA 0.7128 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.995511 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.995511 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.040404 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.040404 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.109989 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.109989 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 6.29 2.29 6.57 2.57 ;
      LAYER ME2 ;
        RECT 6.21 2.21 6.65 2.65 ;
      LAYER ME1 ;
        RECT 8.31 2.2 8.71 2.6 ;
        RECT 6.21 2.31 8.71 2.55 ;
        RECT 6.21 2.23 6.67 2.55 ;
        RECT 6.21 2.23 6.65 2.57 ;
    END
  END CIN
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3712 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2672 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.2156 LAYER ME1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 4.6 3.92 4.88 4.2 ;
        RECT 4.6 1.16 4.88 1.44 ;
      LAYER ME2 ;
        RECT 4.52 3.84 4.96 4.28 ;
        RECT 4.52 1.08 4.96 1.52 ;
        RECT 4.6 1.08 4.88 4.28 ;
      LAYER ME1 ;
        RECT 4.52 1.08 4.96 1.52 ;
        RECT 4.48 1.08 4.96 1.48 ;
        RECT 4.48 3.84 4.96 4.28 ;
        RECT 4.48 3.84 4.88 4.68 ;
    END
  END COUT
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1152 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 11.02 2.02 11.3 2.3 ;
      LAYER ME2 ;
        RECT 10.94 1.94 11.38 2.38 ;
      LAYER ME1 ;
        RECT 10.94 1.94 11.38 2.38 ;
        RECT 10.96 4.06 11.36 4.68 ;
        RECT 11.12 1.08 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
    END
  END S
  OBS
    LAYER ME1 ;
      RECT 0.32 3.36 1.84 3.6 ;
      RECT 1.6 3.36 1.84 4.68 ;
      RECT 0.32 3.36 0.56 4.68 ;
      RECT 0.16 3.84 0.56 4.68 ;
      RECT 1.6 3.84 2 4.68 ;
      RECT 0.16 1.08 0.56 1.48 ;
      RECT 1.6 1.08 2 1.48 ;
      RECT 0.32 1.08 0.56 1.96 ;
      RECT 1.6 1.08 1.84 1.96 ;
      RECT 0.32 1.72 1.84 1.96 ;
      RECT 2.32 3.84 2.76 4.28 ;
      RECT 2.32 3.84 2.72 4.68 ;
      RECT 2.32 1.08 2.72 1.8 ;
      RECT 2.32 1.36 2.76 1.8 ;
      RECT 6.08 3.36 7.6 3.6 ;
      RECT 7.36 3.36 7.6 4.68 ;
      RECT 6.08 3.36 6.32 4.68 ;
      RECT 5.92 3.84 6.32 4.68 ;
      RECT 7.36 3.84 7.76 4.68 ;
      RECT 7.36 1.08 7.84 1.48 ;
      RECT 7.4 1.08 7.84 1.52 ;
      RECT 2.56 2.52 3 2.96 ;
      RECT 3.99 2.56 4.39 2.96 ;
      RECT 2.56 2.72 6.01 2.96 ;
      RECT 5.77 2.88 8.13 3.12 ;
      RECT 7.81 2.84 8.13 3.24 ;
      RECT 8.08 3.48 8.52 3.92 ;
      RECT 8.08 3.48 8.48 4.68 ;
      RECT 8.08 1.08 8.48 1.48 ;
      RECT 9.52 1.08 9.92 1.48 ;
      RECT 8.24 1.08 8.48 1.96 ;
      RECT 9.52 1.08 9.76 1.96 ;
      RECT 8.24 1.72 9.76 1.96 ;
      RECT 8.66 2.96 10.87 3.2 ;
      RECT 8.66 2.84 9.1 3.28 ;
      RECT 10.47 2.88 10.87 3.28 ;
    LAYER ME2 ;
      RECT 2.32 1.36 2.76 1.8 ;
      RECT 2.48 2.52 3 2.96 ;
      RECT 2.48 1.36 2.76 4.28 ;
      RECT 2.32 3.84 2.76 4.28 ;
      RECT 7.4 1.08 7.84 1.52 ;
      RECT 7.56 1.08 7.84 2.28 ;
      RECT 7.56 2 8.52 2.28 ;
      RECT 8.24 2.84 9.1 3.28 ;
      RECT 8.24 2 8.52 3.92 ;
      RECT 8.08 3.48 8.52 3.92 ;
  END
  PROPERTY pathCL "yes" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY instLabel "master" ;
  PROPERTY startLevel 0 ;
  PROPERTY stopLevel 0 ;
  PROPERTY maxDragFig 500 ;
  PROPERTY maxDragLevel 32 ;
  PROPERTY scrollPercent 25 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY instanceDrawingMode "BBox" ;
  PROPERTY lppVisibilityMode "donotCheckValidity" ;
  PROPERTY filterSize 6 ;
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_FA

MACRO UCL_FILL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_FILL 0 0 ;
  SIZE 0.72 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 0.72 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0 4.92 0.72 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 0.72 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0 0.44 0.72 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_FILL

MACRO UCL_GTINVS
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_GTINVS 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.47591 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.47591 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.076696 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.076696 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.192724 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.192724 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
    END
  END EN
  PIN AUS
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 2.74 2.66 3.02 ;
      LAYER ME2 ;
        RECT 2.3 2.66 2.74 3.1 ;
      LAYER ME1 ;
        RECT 2.3 2.66 2.74 3.1 ;
        RECT 2.32 3.56 2.72 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 2.43 1.08 2.67 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2616 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.798535 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.798535 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.02 1.94 2.3 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.02 2.38 ;
      LAYER ME1 ;
        RECT 1.58 1.96 2.19 2.36 ;
        RECT 1.58 1.94 2.02 2.38 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.16 1.08 0.56 1.48 ;
      RECT 1.07 2.8 1.47 3.2 ;
      RECT 0.24 2.96 1.47 3.2 ;
      RECT 0.24 1.08 0.48 4.68 ;
      RECT 0.16 3.56 0.56 4.68 ;
      RECT 1.6 3.56 2 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_GTINVS

MACRO UCL_ICG
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_ICG 0 0 ;
  SIZE 12.24 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 3.74 2.67 4.18 3.11 ;
        RECT 3.74 2.69 4.39 3.09 ;
    END
  END EN
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.94 1.94 11.38 2.38 ;
    END
  END GCLK
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 12.24 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.76 0.44 4.16 1.48 ;
        RECT 6.64 0.44 7.04 1.48 ;
        RECT 8.08 0.44 8.48 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 0 0.44 12.24 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 12.24 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.76 3.56 4.16 5.32 ;
        RECT 6.64 3.56 7.04 5.32 ;
        RECT 8.08 3.56 8.48 5.32 ;
        RECT 9.52 3.56 9.92 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 0 4.92 12.24 5.32 ;
    END
  END vddd
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3824 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.1568 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.343101 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.343101 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.21978 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.21978 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.478632 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.478632 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.92 0.5 3.2 ;
        RECT 0.22 2.36 0.5 2.64 ;
        RECT 8.14 2.02 8.42 2.3 ;
      LAYER ME1 ;
        RECT 8.06 1.94 8.5 2.38 ;
        RECT 0.14 2.28 0.58 3.28 ;
      LAYER ME2 ;
        RECT 8.06 1.94 8.5 2.38 ;
        RECT 0.22 2.02 8.5 2.3 ;
        RECT 0.22 2.02 0.5 3.28 ;
    END
  END CLK
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 2.04 2.06 2.28 ;
      RECT 1.58 1.97 2.06 2.37 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 1.58 1.95 2.02 2.39 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 2.4 1.76 2.91 2.16 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 3.04 1.08 3.44 1.48 ;
      RECT 3.2 2.19 5.11 2.43 ;
      RECT 4.71 2.19 5.11 2.59 ;
      RECT 3.2 1.08 3.44 4.68 ;
      RECT 3.04 3.56 3.44 4.68 ;
      RECT 5.2 1.08 5.6 1.48 ;
      RECT 5.36 2.77 7.23 3.01 ;
      RECT 6.83 2.69 7.23 3.09 ;
      RECT 5.36 1.08 5.6 4.68 ;
      RECT 5.2 3.56 5.6 4.68 ;
      RECT 7.36 1.08 7.76 1.48 ;
      RECT 6.22 2.05 7.78 2.29 ;
      RECT 6.22 1.96 6.62 2.36 ;
      RECT 9.03 1.96 9.43 2.36 ;
      RECT 7.34 1.95 7.78 2.39 ;
      RECT 9.03 1.96 9.36 2.45 ;
      RECT 8.82 2.44 9.27 2.57 ;
      RECT 8.94 2.35 9.03 2.78 ;
      RECT 8.72 2.56 9.15 2.69 ;
      RECT 8.06 2.66 9.03 2.78 ;
      RECT 7.47 2.76 8.94 2.9 ;
      RECT 7.47 2.76 8.5 3 ;
      RECT 8.06 2.66 8.5 3.1 ;
      RECT 7.47 1.08 7.71 4.68 ;
      RECT 7.36 3.56 7.76 4.68 ;
      RECT 9.52 1.08 9.92 1.48 ;
      RECT 9.68 1.08 9.92 3.1 ;
      RECT 9.32 2.82 9.44 3.28 ;
      RECT 9.2 2.94 10.66 3.1 ;
      RECT 9.44 2.76 9.5 3.16 ;
      RECT 9.16 3.06 10.66 3.1 ;
      RECT 9.5 2.66 10.66 3.1 ;
      RECT 9.04 3.1 9.44 3.28 ;
      RECT 8.92 3.22 9.32 3.4 ;
      RECT 8.8 3.34 9.2 4.68 ;
  END
END UCL_ICG

MACRO UCL_INV
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV

MACRO UCL_INV16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV16 0 0 ;
  SIZE 30.24 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 5.92 3.56 6.32 5.32 ;
        RECT 7.36 3.56 7.76 5.32 ;
        RECT 8.8 3.56 9.2 5.32 ;
        RECT 10.24 3.56 10.64 5.32 ;
        RECT 11.68 3.56 12.08 5.32 ;
        RECT 13.12 3.56 13.52 5.32 ;
        RECT 14.56 3.56 14.96 5.32 ;
        RECT 16 3.56 16.4 5.32 ;
        RECT 17.44 3.56 17.84 5.32 ;
        RECT 18.88 3.56 19.28 5.32 ;
        RECT 20.32 3.56 20.72 5.32 ;
        RECT 21.76 3.56 22.16 5.32 ;
        RECT 23.2 3.56 23.6 5.32 ;
        RECT 24.64 3.56 25.04 5.32 ;
        RECT 26.08 3.56 26.48 5.32 ;
        RECT 27.52 3.56 27.92 5.32 ;
        RECT 28.96 3.56 29.36 5.32 ;
        RECT 0 4.92 30.24 5.32 ;
    END
  END vddd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.7232 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 75.0336 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 1.2544 LAYER VI1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME1 ;
    ANTENNADIFFAREA 14.2688 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 8.14 2.02 8.42 2.3 ;
        RECT 9.58 2.02 9.86 2.3 ;
        RECT 11.02 2.02 11.3 2.3 ;
        RECT 12.46 2.02 12.74 2.3 ;
        RECT 13.9 2.02 14.18 2.3 ;
        RECT 15.34 2.02 15.62 2.3 ;
        RECT 16.78 2.02 17.06 2.3 ;
        RECT 18.22 2.02 18.5 2.3 ;
        RECT 19.66 2.02 19.94 2.3 ;
        RECT 21.1 2.02 21.38 2.3 ;
        RECT 22.54 2.02 22.82 2.3 ;
        RECT 23.98 2.02 24.26 2.3 ;
        RECT 25.42 2.02 25.7 2.3 ;
        RECT 26.86 2.02 27.14 2.3 ;
        RECT 28.3 2.02 28.58 2.3 ;
        RECT 29.74 2.02 30.02 2.3 ;
      LAYER ME2 ;
        RECT 8.06 1.94 30.1 2.38 ;
      LAYER ME1 ;
        RECT 8.06 1.94 30.1 2.38 ;
        RECT 29.68 3.56 30.08 4.68 ;
        RECT 29.68 1.08 30.08 1.48 ;
        RECT 29.76 1.08 30 4.68 ;
        RECT 28.24 3.56 28.64 4.68 ;
        RECT 28.24 1.08 28.64 1.48 ;
        RECT 28.32 1.08 28.56 4.68 ;
        RECT 26.8 3.56 27.2 4.68 ;
        RECT 26.8 1.08 27.2 1.48 ;
        RECT 26.88 1.08 27.12 4.68 ;
        RECT 25.36 3.56 25.76 4.68 ;
        RECT 25.36 1.08 25.76 1.48 ;
        RECT 25.44 1.08 25.68 4.68 ;
        RECT 23.92 3.56 24.32 4.68 ;
        RECT 23.92 1.08 24.32 1.48 ;
        RECT 24 1.08 24.24 4.68 ;
        RECT 22.48 3.56 22.88 4.68 ;
        RECT 22.48 1.08 22.88 1.48 ;
        RECT 22.56 1.08 22.8 4.68 ;
        RECT 21.04 3.56 21.44 4.68 ;
        RECT 21.04 1.08 21.44 1.48 ;
        RECT 21.12 1.08 21.36 4.68 ;
        RECT 19.6 3.56 20 4.68 ;
        RECT 19.6 1.08 20 1.48 ;
        RECT 19.68 1.08 19.92 4.68 ;
        RECT 18.16 3.56 18.56 4.68 ;
        RECT 18.16 1.08 18.56 1.48 ;
        RECT 18.24 1.08 18.48 4.68 ;
        RECT 16.72 3.56 17.12 4.68 ;
        RECT 16.72 1.08 17.12 1.48 ;
        RECT 16.8 1.08 17.04 4.68 ;
        RECT 15.28 3.56 15.68 4.68 ;
        RECT 15.28 1.08 15.68 1.48 ;
        RECT 15.36 1.08 15.6 4.68 ;
        RECT 13.84 3.56 14.24 4.68 ;
        RECT 13.84 1.08 14.24 1.48 ;
        RECT 13.92 1.08 14.16 4.68 ;
        RECT 12.4 3.56 12.8 4.68 ;
        RECT 12.4 1.08 12.8 1.48 ;
        RECT 12.48 1.08 12.72 4.68 ;
        RECT 10.96 3.56 11.36 4.68 ;
        RECT 10.96 1.08 11.36 1.48 ;
        RECT 11.04 1.08 11.28 4.68 ;
        RECT 9.52 3.56 9.92 4.68 ;
        RECT 9.52 1.08 9.92 1.48 ;
        RECT 9.6 1.08 9.84 4.68 ;
        RECT 8.08 3.56 8.48 4.68 ;
        RECT 8.08 1.08 8.48 1.48 ;
        RECT 8.16 1.08 8.4 4.68 ;
    END
  END AUS
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 5.92 0.44 6.32 1.48 ;
        RECT 7.36 0.44 7.76 1.48 ;
        RECT 8.8 0.44 9.2 1.48 ;
        RECT 10.24 0.44 10.64 1.48 ;
        RECT 11.68 0.44 12.08 1.48 ;
        RECT 13.12 0.44 13.52 1.48 ;
        RECT 14.56 0.44 14.96 1.48 ;
        RECT 16 0.44 16.4 1.48 ;
        RECT 17.44 0.44 17.84 1.48 ;
        RECT 18.88 0.44 19.28 1.48 ;
        RECT 20.32 0.44 20.72 1.48 ;
        RECT 21.76 0.44 22.16 1.48 ;
        RECT 23.2 0.44 23.6 1.48 ;
        RECT 24.64 0.44 25.04 1.48 ;
        RECT 26.08 0.44 26.48 1.48 ;
        RECT 27.52 0.44 27.92 1.48 ;
        RECT 28.96 0.44 29.36 1.48 ;
        RECT 0 0.44 30.24 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 30.24 5.96 ;
    END
  END vddb
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 30.24 0.2 ;
    END
  END gndb
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.86 1.94 1.3 2.38 ;
      RECT 0.96 2.66 2.02 3.1 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 3.02 2.66 3.46 3.1 ;
      RECT 4.46 2.66 4.9 3.1 ;
      RECT 5.9 2.66 6.34 3.1 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 5.2 1.08 5.6 1.48 ;
      RECT 6.64 1.08 7.04 1.48 ;
      RECT 2.3 1.94 7.26 2.38 ;
      RECT 6.72 1.94 7.26 3.1 ;
      RECT 6.72 2.66 7.78 3.1 ;
      RECT 2.4 1.08 2.64 4.68 ;
      RECT 3.84 1.08 4.08 4.68 ;
      RECT 5.28 1.08 5.52 4.68 ;
      RECT 6.72 1.08 6.96 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
      RECT 5.2 3.56 5.6 4.68 ;
      RECT 6.64 3.56 7.04 4.68 ;
      RECT 8.78 2.66 9.22 3.1 ;
      RECT 10.22 2.66 10.66 3.1 ;
      RECT 11.66 2.66 12.1 3.1 ;
      RECT 13.1 2.66 13.54 3.1 ;
      RECT 14.54 2.66 14.98 3.1 ;
      RECT 15.98 2.66 16.42 3.1 ;
      RECT 17.42 2.66 17.86 3.1 ;
      RECT 18.86 2.66 19.3 3.1 ;
      RECT 20.3 2.66 20.74 3.1 ;
      RECT 21.74 2.66 22.18 3.1 ;
      RECT 23.18 2.66 23.62 3.1 ;
      RECT 24.62 2.66 25.06 3.1 ;
      RECT 26.06 2.66 26.5 3.1 ;
      RECT 27.5 2.66 27.94 3.1 ;
      RECT 28.94 2.66 29.38 3.1 ;
    LAYER ME2 ;
      RECT 6.72 2.66 29.38 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV16

MACRO UCL_INV2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV2 0 0 ;
  SIZE 2.16 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.16 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 0 4.92 2.16 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.16 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 2.16 0.84 ;
    END
  END gndd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.96 1.08 1.2 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 0.86 1.94 1.3 2.38 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV2

MACRO UCL_INV4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV4 0 0 ;
  SIZE 5.76 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1008 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3552 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 3.5672 LAYER ME1 ;
    ANTENNADIFFAREA 3.5672 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 5.26 2.02 5.54 2.3 ;
      LAYER ME2 ;
        RECT 5.18 1.94 5.62 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 5.62 2.38 ;
        RECT 5.2 3.56 5.6 4.68 ;
        RECT 5.2 1.08 5.6 1.48 ;
        RECT 5.28 1.08 5.52 4.68 ;
        RECT 3.76 3.56 4.16 4.68 ;
        RECT 3.76 1.08 4.16 1.48 ;
        RECT 3.84 1.08 4.08 4.68 ;
        RECT 2.32 3.56 2.72 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 2.4 1.08 2.64 4.68 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7744 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.3792 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.3104 LAYER ME1 ;
      ANTENNAGATEAREA 1.3104 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.059829 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.059829 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 5.76 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 0 4.92 5.76 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 5.76 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 0 0.44 5.76 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 1.58 2.66 2.02 3.1 ;
      RECT 3.02 2.66 3.46 3.1 ;
      RECT 4.46 2.66 4.9 3.1 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV4

MACRO UCL_INV_LP
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV_LP 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME1 ;
    ANTENNADIFFAREA 0.4312 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
        RECT 0.88 4.28 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME1 ;
      ANTENNAGATEAREA 0.1584 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.222222 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.222222 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.333333 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.333333 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.494949 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 4.28 0.56 5.32 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV_LP

MACRO UCL_INV_LP2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_INV_LP2 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1152 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME1 ;
    ANTENNADIFFAREA 0.6468 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
        RECT 0.88 4.06 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.814815 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.814815 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.555556 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.555556 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 4.06 0.56 5.32 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_INV_LP2

MACRO UCL_LAT
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_LAT 0 0 ;
  SIZE 6.48 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.3 2.67 2.74 3.11 ;
        RECT 2.3 2.69 2.95 3.09 ;
    END
  END A
  PIN L
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.95 0.58 2.39 ;
        RECT 0.14 1.97 0.62 2.37 ;
    END
  END L
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 4.78 1.96 5.18 2.36 ;
        RECT 4.78 2.05 6.34 2.29 ;
        RECT 6.03 1.08 6.27 4.68 ;
        RECT 5.92 1.08 6.32 1.48 ;
        RECT 5.92 3.56 6.32 4.68 ;
        RECT 5.9 1.95 6.34 2.39 ;
    END
  END Q
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 6.48 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.32 0.44 2.72 1.48 ;
        RECT 5.2 0.44 5.6 1.48 ;
        RECT 0 0.44 6.48 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 6.48 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 5.2 3.56 5.6 5.32 ;
        RECT 0 4.92 6.48 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.96 1.76 1.47 2.16 ;
      RECT 0.96 1.08 1.2 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 1.6 1.08 2 1.48 ;
      RECT 1.76 2.19 3.67 2.43 ;
      RECT 3.27 2.19 3.67 2.59 ;
      RECT 1.76 1.08 2 4.68 ;
      RECT 1.6 3.56 2 4.68 ;
      RECT 3.76 1.08 4.16 1.48 ;
      RECT 3.92 2.77 5.79 3.01 ;
      RECT 5.39 2.69 5.79 3.09 ;
      RECT 3.92 1.08 4.16 4.68 ;
      RECT 3.76 3.56 4.16 4.68 ;
  END
END UCL_LAT

MACRO UCL_MUX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_MUX2 0 0 ;
  SIZE 4.32 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0464 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.79 3.1 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27365 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.438528 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9828 LAYER ME1 ;
    ANTENNADIFFAREA 0.9828 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 1.34 3.56 1.74 4.68 ;
        RECT 1.34 1.08 1.74 1.48 ;
        RECT 1.25 3.49 1.65 3.58 ;
        RECT 1.21 3.37 1.58 3.5 ;
        RECT 1.34 1.08 1.58 2.07 ;
        RECT 1.09 3.25 1.46 3.46 ;
        RECT 0.86 1.94 1.46 2.19 ;
        RECT 1.09 3.24 1.34 3.46 ;
        RECT 1.33 3.56 1.74 3.59 ;
        RECT 1.25 1.86 1.58 2.07 ;
        RECT 1.33 1.85 1.34 2.2 ;
        RECT 1.09 1.94 1.33 3.46 ;
        RECT 0.86 1.94 1.33 2.38 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3124 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.104 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 2.02 2.66 2.3 ;
      LAYER ME2 ;
        RECT 2.3 1.94 2.74 2.38 ;
      LAYER ME1 ;
        RECT 2.03 1.94 2.74 2.38 ;
    END
  END EIN0
  PIN SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1484 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.928 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.82 2.74 4.1 3.02 ;
      LAYER ME2 ;
        RECT 3.74 2.66 4.18 3.1 ;
      LAYER ME1 ;
        RECT 1.57 2.66 4.18 3.1 ;
    END
  END SEL
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 4.32 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 2.52 3.56 2.92 5.32 ;
        RECT 0 4.92 4.32 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 4.32 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 2.52 0.44 2.92 1.48 ;
        RECT 0 0.44 4.32 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 3.24 3.56 4.18 4.46 ;
      RECT 3.24 3.56 3.64 4.68 ;
      RECT 3.24 1.08 4.18 1.48 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_MUX2

MACRO UCL_MUX2A
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_MUX2A 0 0 ;
  SIZE 5.04 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0464 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.873016 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.74 1.22 3.02 ;
      LAYER ME2 ;
        RECT 0.86 2.66 1.3 3.1 ;
      LAYER ME1 ;
        RECT 0.65 2.66 1.3 3.1 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30045 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.528505 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9828 LAYER ME1 ;
    ANTENNADIFFAREA 0.9828 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 3.46 1.94 3.74 ;
      LAYER ME2 ;
        RECT 1.58 3.38 2.02 3.82 ;
      LAYER ME1 ;
        RECT 2.06 3.56 2.46 4.68 ;
        RECT 2.06 1.08 2.46 1.48 ;
        RECT 2.06 1.08 2.3 2.07 ;
        RECT 1.81 1.98 2.18 2.19 ;
        RECT 1.58 3.52 2.1 3.82 ;
        RECT 1.58 3.51 2.06 3.82 ;
        RECT 2.05 3.56 2.46 3.86 ;
        RECT 1.93 1.89 2.3 2.07 ;
        RECT 2.05 1.85 2.06 2.2 ;
        RECT 1.58 3.38 2.05 3.82 ;
        RECT 1.81 1.98 2.05 3.82 ;
        RECT 2.02 1.86 2.05 3.85 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3124 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.104 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.953602 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.369963 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 3.1 2.02 3.38 2.3 ;
      LAYER ME2 ;
        RECT 3.02 1.94 3.46 2.38 ;
      LAYER ME1 ;
        RECT 2.75 1.94 3.46 2.38 ;
    END
  END EIN0
  PIN SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1484 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.928 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.752747 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 4.468864 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 4.54 2.74 4.82 3.02 ;
      LAYER ME2 ;
        RECT 4.46 2.66 4.9 3.1 ;
      LAYER ME1 ;
        RECT 2.29 2.66 4.9 3.1 ;
    END
  END SEL
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 5.04 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 3.24 3.56 3.64 5.32 ;
        RECT 0 4.92 5.04 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 5.04 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 3.24 0.44 3.64 1.48 ;
        RECT 0 0.44 5.04 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.16 1.08 0.56 1.48 ;
      RECT 0.16 1.81 1.51 2.05 ;
      RECT 1.11 1.73 1.51 2.13 ;
      RECT 0.16 1.08 0.4 4.68 ;
      RECT 0.16 3.56 0.56 4.68 ;
      RECT 3.96 3.56 4.9 4.46 ;
      RECT 3.96 3.56 4.36 4.68 ;
      RECT 3.96 1.08 4.9 1.48 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_MUX2A

MACRO UCL_MUX2B
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_MUX2B 0 0 ;
  SIZE 5.04 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 5.04 5.96 ;
    END
  END vddb
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 5.04 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 3.24 0.44 3.64 1.48 ;
        RECT 0 0.44 5.04 0.84 ;
    END
  END gndd
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 3.24 3.56 3.64 5.32 ;
        RECT 0 4.92 5.04 5.32 ;
    END
  END vddd
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.11 1.73 1.51 2.18 ;
    END
  END EIN1
  PIN SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.29 2.66 4.9 3.1 ;
    END
  END SEL
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.16 1.08 0.4 4.68 ;
        RECT 0.16 1.08 0.56 1.48 ;
        RECT 0.16 3.56 0.56 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.75 1.94 3.46 2.38 ;
    END
  END EIN0
  OBS
    LAYER ME1 ;
      RECT 2.06 1.08 2.46 1.48 ;
      RECT 2.05 1.85 2.06 2.2 ;
      RECT 2.06 1.08 2.3 2.07 ;
      RECT 1.81 1.98 2.18 2.19 ;
      RECT 0.65 2.76 2.05 3 ;
      RECT 0.65 2.68 1.05 3.08 ;
      RECT 1.81 3.52 2.1 3.73 ;
      RECT 1.81 1.98 2.05 3.73 ;
      RECT 1.93 1.86 2.05 3.85 ;
      RECT 2.05 3.51 2.06 3.86 ;
      RECT 2.06 3.56 2.46 4.68 ;
      RECT 3.96 3.56 4.9 4.46 ;
      RECT 3.96 3.56 4.36 4.68 ;
      RECT 3.96 1.08 4.9 1.48 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_MUX2B

MACRO UCL_NAND2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NAND2 0 0 ;
  SIZE 2.16 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5096 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.824 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.555556 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.555556 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.567766 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.567766 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.1 1.96 1.5 2.36 ;
        RECT 0.14 2.01 1.5 2.31 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3736 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6848 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9608 LAYER ME1 ;
    ANTENNADIFFAREA 0.9608 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.74 1.94 3.02 ;
      LAYER ME2 ;
        RECT 1.58 2.66 2.02 3.1 ;
      LAYER ME1 ;
        RECT 1.02 2.84 2.02 3.1 ;
        RECT 1.58 2.66 2.02 3.1 ;
        RECT 1.74 1.08 2 3.1 ;
        RECT 1.6 1.08 2 1.48 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 1.02 2.84 1.28 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.590965 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.578755 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.16 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 0 4.92 2.16 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.16 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 2.16 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NAND2

MACRO UCL_NAND2A
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NAND2A 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2496 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9792 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.761905 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.761905 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.989011 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.989011 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.74 1.22 3.02 ;
      LAYER ME2 ;
        RECT 0.86 2.66 1.3 3.1 ;
      LAYER ME1 ;
        RECT 0.86 2.66 1.3 3.1 ;
        RECT 0.72 2.69 1.3 3.09 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4888 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.704 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9608 LAYER ME1 ;
    ANTENNADIFFAREA 0.9608 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 1.3 2.66 1.58 ;
      LAYER ME2 ;
        RECT 2.3 1.22 2.74 1.66 ;
      LAYER ME1 ;
        RECT 1.6 2.88 2.74 3.12 ;
        RECT 2.46 1.22 2.74 3.12 ;
        RECT 2.32 1.08 2.72 1.66 ;
        RECT 2.3 1.22 2.74 1.66 ;
        RECT 1.6 2.88 2 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2256 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9216 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.688645 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.688645 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.813187 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.813187 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.75 2.02 2.03 2.3 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.11 2.38 ;
      LAYER ME1 ;
        RECT 1.67 1.96 2.19 2.36 ;
        RECT 1.67 1.94 2.11 2.38 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.88 3.56 1.28 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.88 0.44 1.28 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.16 1.08 0.56 1.48 ;
      RECT 0.24 1.91 1.43 2.15 ;
      RECT 1.11 1.83 1.43 2.23 ;
      RECT 0.24 1.08 0.48 4.68 ;
      RECT 0.16 3.56 0.56 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NAND2A

MACRO UCL_NAND2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NAND2_2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 3.04 0.44 3.44 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8136 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.13 2.06 2.71 2.46 ;
        RECT 2.3 1.94 2.74 2.38 ;
    END
  END EIN1
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9656 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.02 2.84 1.28 4.68 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 1.6 1.08 1.86 3.1 ;
        RECT 1.6 1.08 2 1.66 ;
        RECT 1.58 1.22 2.02 1.66 ;
        RECT 1.02 2.84 2.58 3.1 ;
        RECT 2.32 2.84 2.58 4.68 ;
        RECT 2.32 3.56 2.72 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8136 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NAND2_2

MACRO UCL_NAND2_WIDEN
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NAND2_WIDEN 0 0 ;
  SIZE 2.16 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 0 4.92 2.16 5.32 ;
    END
  END vddd
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 2.16 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.16 5.96 ;
    END
  END vddb
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.46 ;
        RECT 0.85 2.06 1.44 2.46 ;
    END
  END EIN1
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.16 0.2 ;
    END
  END gndb
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1764 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.02 2.84 1.28 4.68 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 1.6 1.08 2 1.48 ;
        RECT 1.74 1.08 2 3.1 ;
        RECT 1.58 2.66 2.02 3.1 ;
        RECT 1.02 2.84 2.02 3.1 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NAND2_WIDEN

MACRO UCL_NAND3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NAND3 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.84 0.56 5.32 ;
        RECT 1.6 3.84 2 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.46 ;
        RECT 0.85 2.06 1.44 2.46 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.58 1.22 2.02 1.66 ;
        RECT 1.78 1.22 2.02 2.46 ;
        RECT 1.78 2.06 2.19 2.46 ;
    END
  END EIN2
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3376 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.02 2.84 1.28 4.68 ;
        RECT 0.88 3.84 1.28 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 1.02 2.84 2.72 3.1 ;
        RECT 2.46 1.08 2.72 4.68 ;
        RECT 2.32 3.38 2.72 4.68 ;
        RECT 2.3 3.38 2.74 3.82 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3168 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NAND3

MACRO UCL_NOR2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NOR2 0 0 ;
  SIZE 2.16 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.111552 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.742268 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.742268 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 6.046827 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 6.046827 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.11 2.68 1.51 3.08 ;
        RECT 1.03 2.59 1.44 2.7 ;
        RECT 0.91 2.47 1.35 2.62 ;
        RECT 0.79 2.35 1.23 2.5 ;
        RECT 0.14 2.27 1.11 2.38 ;
        RECT 0.14 2.15 1.03 2.38 ;
        RECT 0.14 2.03 0.91 2.38 ;
        RECT 0.14 1.94 0.79 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2834 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.467811 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9726 LAYER ME1 ;
    ANTENNADIFFAREA 0.9726 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.02 1.94 2.3 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.02 2.38 ;
      LAYER ME1 ;
        RECT 1.58 1.94 2.02 2.38 ;
        RECT 1.6 3.56 2 4.68 ;
        RECT 1.76 1.94 2 4.68 ;
        RECT 1.16 1.88 1.58 1.99 ;
        RECT 1.52 1.94 2.02 2.29 ;
        RECT 1.16 1.76 1.52 1.99 ;
        RECT 1.4 1.94 2.02 2.23 ;
        RECT 1.04 1.64 1.4 1.87 ;
        RECT 1.28 1.94 2.02 2.11 ;
        RECT 1.04 1.08 1.28 1.87 ;
        RECT 0.88 1.08 1.28 1.48 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.16 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 0 4.92 2.16 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.16 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 2.16 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NOR2

MACRO UCL_NOR2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NOR2_2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.111552 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.928571 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.928571 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.222759 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.222759 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.11 2.68 1.51 3.08 ;
        RECT 1.03 2.59 1.44 2.7 ;
        RECT 0.91 2.47 1.35 2.62 ;
        RECT 0.79 2.35 1.23 2.5 ;
        RECT 0.14 2.27 1.11 2.38 ;
        RECT 0.14 2.15 1.03 2.38 ;
        RECT 0.14 2.03 0.91 2.38 ;
        RECT 0.14 1.94 0.79 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2834 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.467811 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 1.2204 LAYER ME1 ;
    ANTENNADIFFAREA 1.2204 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.02 1.94 2.3 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.02 2.38 ;
      LAYER ME1 ;
        RECT 1.58 1.94 2.02 2.38 ;
        RECT 1.6 3.56 2 4.68 ;
        RECT 1.76 1.94 2 4.68 ;
        RECT 1.16 1.88 1.58 1.99 ;
        RECT 1.52 1.94 2.02 2.29 ;
        RECT 1.16 1.76 1.52 1.99 ;
        RECT 1.4 1.94 2.02 2.23 ;
        RECT 1.04 1.64 1.4 1.87 ;
        RECT 1.28 1.94 2.02 2.11 ;
        RECT 1.04 1.08 1.28 1.87 ;
        RECT 0.88 1.08 1.28 1.48 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.295482 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.295482 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 1.289377 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 1.289377 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 3.04 3.56 3.44 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NOR2_2

MACRO UCL_NOR3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_NOR3 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.86 2.66 1.3 3.1 ;
        RECT 0.86 2.68 1.47 3.08 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.78 2.76 2.02 3.82 ;
        RECT 1.58 3.38 2.02 3.82 ;
        RECT 1.78 2.76 2.15 3.16 ;
    END
  END EIN2
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.345 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 1.04 1.08 1.28 1.96 ;
        RECT 1.04 1.72 2.63 1.96 ;
        RECT 2.39 1.08 2.63 4.68 ;
        RECT 2.32 1.08 2.72 1.48 ;
        RECT 2.32 3.56 2.72 4.68 ;
        RECT 2.3 4.1 2.74 4.54 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4068 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN0
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_NOR3

MACRO UCL_OAI21
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_OAI21 0 0 ;
  SIZE 2.88 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 2.88 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 0 0.44 2.88 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 2.88 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 4.06 0.56 5.32 ;
        RECT 2.32 4.06 2.72 5.32 ;
        RECT 0 4.92 2.88 5.32 ;
    END
  END vddd
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1792 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.5696 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.9108 LAYER ME1 ;
    ANTENNADIFFAREA 0.9108 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 4.18 1.22 4.46 ;
      LAYER ME2 ;
        RECT 0.86 4.1 1.3 4.54 ;
      LAYER ME1 ;
        RECT 0.86 4.1 1.3 4.54 ;
        RECT 0.88 4.06 1.28 4.68 ;
        RECT 0.88 2.2 1.12 4.68 ;
        RECT 0.32 2.2 1.12 2.44 ;
        RECT 0.32 1.08 0.56 2.44 ;
        RECT 0.16 1.08 0.56 1.48 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2056 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8736 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.627595 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.627595 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.666667 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.666667 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 2.38 2.28 2.66 2.56 ;
      LAYER ME2 ;
        RECT 2.3 1.94 2.74 2.64 ;
      LAYER ME1 ;
        RECT 2.3 2.2 2.74 2.64 ;
        RECT 2.27 2.22 2.74 2.62 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2776 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0464 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.847375 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.847375 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.194139 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.239316 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.74 1.94 3.02 ;
      LAYER ME2 ;
        RECT 1.58 2.66 2.02 3.1 ;
      LAYER ME1 ;
        RECT 1.58 2.66 2.02 3.1 ;
        RECT 1.37 2.68 2.02 3.08 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1968 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8544 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME1 ;
      ANTENNAGATEAREA 0.2376 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.828283 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.828283 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 3.59596 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 3.59596 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.329966 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.68 0.61 3.08 ;
        RECT 0.14 2.68 0.58 3.1 ;
    END
  END EIN2
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 1.04 1.08 1.28 1.96 ;
      RECT 2.32 1.08 2.56 1.96 ;
      RECT 1.04 1.72 2.56 1.96 ;
  END
END UCL_OAI21

MACRO UCL_OAI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_OAI22 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2326 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.95 1.81 1.19 4.54 ;
        RECT 0.86 4.1 1.3 4.54 ;
        RECT 0.95 1.81 1.35 2.21 ;
        RECT 0.95 4.06 2 4.3 ;
        RECT 1.6 4.06 2 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.89 1.96 3.46 2.36 ;
        RECT 3.02 1.94 3.46 2.38 ;
    END
  END EIN0
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 2.2 2.68 2.74 3.08 ;
        RECT 2.3 2.66 2.74 3.1 ;
    END
  END EIN1
  PIN EIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
        RECT 0.14 1.96 0.71 2.36 ;
    END
  END EIN2
  PIN EIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3276 LAYER ME1 ;
    PORT
      LAYER ME1 ;
        RECT 1.43 2.68 1.67 3.82 ;
        RECT 1.43 3.38 2.02 3.82 ;
    END
  END EIN3
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 2.25 0.44 2.65 1.08 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 4.06 0.56 5.32 ;
        RECT 3.04 4.06 3.44 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  OBS
    LAYER ME1 ;
      RECT 0.16 1.08 0.56 1.56 ;
      RECT 1.53 1.11 1.93 1.56 ;
      RECT 3.04 1.08 3.44 1.56 ;
      RECT 0.16 1.32 3.44 1.56 ;
  END
END UCL_OAI22

MACRO UCL_OR2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_OR2 0 0 ;
  SIZE 3.6 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.111552 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.742268 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.742268 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 6.046827 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 6.046827 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 1.11 2.68 1.51 3.08 ;
        RECT 1.03 2.59 1.44 2.7 ;
        RECT 0.91 2.47 1.35 2.62 ;
        RECT 0.79 2.35 1.23 2.5 ;
        RECT 0.14 2.27 1.11 2.38 ;
        RECT 0.14 2.15 1.03 2.38 ;
        RECT 0.14 2.03 0.91 2.38 ;
        RECT 0.14 1.94 0.79 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 3.1 2.02 3.38 2.3 ;
      LAYER ME2 ;
        RECT 3.02 1.94 3.46 2.38 ;
      LAYER ME1 ;
        RECT 3.02 1.94 3.46 2.38 ;
        RECT 3.04 3.56 3.44 4.68 ;
        RECT 3.04 1.08 3.44 1.48 ;
        RECT 3.12 1.08 3.36 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME1 ;
      ANTENNAGATEAREA 0.3492 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.55441 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 2.419244 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.224513 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.74 0.5 3.02 ;
      LAYER ME2 ;
        RECT 0.14 2.66 0.58 3.1 ;
      LAYER ME1 ;
        RECT 0.14 2.66 0.58 3.1 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 3.6 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 2.32 3.56 2.72 5.32 ;
        RECT 0 4.92 3.6 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 3.6 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 2.32 0.44 2.72 1.48 ;
        RECT 0 0.44 3.6 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 1.04 1.08 1.28 1.87 ;
      RECT 1.16 1.08 1.28 1.99 ;
      RECT 1.28 1.64 1.4 2.11 ;
      RECT 1.4 1.76 1.52 2.23 ;
      RECT 1.52 1.88 1.58 2.29 ;
      RECT 1.58 1.94 2.02 2.38 ;
      RECT 1.76 2.66 2.74 3.1 ;
      RECT 1.76 1.94 2 4.68 ;
      RECT 1.6 3.56 2 4.68 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_OR2

MACRO UCL_TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_TIEHI 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0.32 0.44 0.56 3.08 ;
        RECT 0.16 2.68 0.56 3.08 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.64 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
END UCL_TIEHI

MACRO UCL_TIELOW
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_TIELOW 0 0 ;
  SIZE 1.44 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1952 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1856 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME1 ;
    ANTENNADIFFAREA 0.8918 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 0.94 2.02 1.22 2.3 ;
      LAYER ME2 ;
        RECT 0.86 1.94 1.3 2.38 ;
      LAYER ME1 ;
        RECT 0.86 1.94 1.3 2.38 ;
        RECT 0.88 3.56 1.28 4.68 ;
        RECT 0.88 1.08 1.28 1.48 ;
        RECT 0.96 1.08 1.2 4.68 ;
    END
  END AUS
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 1.44 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 0.16 2.68 0.56 3.08 ;
        RECT 0.32 2.68 0.56 5.32 ;
        RECT 0.16 3.56 0.56 5.32 ;
        RECT 0 4.92 1.44 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 1.44 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 0.16 0.44 0.56 1.48 ;
        RECT 0 0.44 1.44 0.84 ;
    END
  END gndd
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 0 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_TIELOW

MACRO UCL_XOR
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN UCL_XOR 0 0 ;
  SIZE 6.48 BY 5.76 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN EIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1936 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8448 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 0.295482 LAYER ME1 ;
      ANTENNAMAXAREACAR 0.295482 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 1.289377 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 1.289377 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 0.22 2.02 0.5 2.3 ;
      LAYER ME2 ;
        RECT 0.14 1.94 0.58 2.38 ;
      LAYER ME1 ;
        RECT 0.14 1.94 0.58 2.38 ;
    END
  END EIN1
  PIN AUS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.95 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 10.538539 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNADIFFAREA 1.7836 LAYER ME1 ;
    ANTENNADIFFAREA 1.7836 LAYER ME2 ;
    PORT
      LAYER VI1 ;
        RECT 5.98 1.3 6.26 1.58 ;
      LAYER ME2 ;
        RECT 5.9 1.22 6.34 1.66 ;
      LAYER ME1 ;
        RECT 5.9 1.22 6.34 1.66 ;
        RECT 5.92 3.56 6.32 4.68 ;
        RECT 5.9 1.08 6.32 1.66 ;
        RECT 5.99 1.08 6.23 4.68 ;
        RECT 5.45 1.24 6.34 1.48 ;
        RECT 5.09 1.5 5.47 1.6 ;
        RECT 4.99 1.62 5.45 1.72 ;
        RECT 5.09 1.5 5.45 1.72 ;
        RECT 5.21 1.38 5.57 1.58 ;
        RECT 5.33 1.26 5.45 1.72 ;
        RECT 4.14 1.72 5.33 1.84 ;
        RECT 4.26 1.72 5.21 1.96 ;
        RECT 4.02 1.62 4.38 1.82 ;
        RECT 3.9 1.6 4.28 1.7 ;
        RECT 3.9 1.48 4.26 1.7 ;
        RECT 4.14 1.72 5.21 1.94 ;
        RECT 3.04 1.36 4.14 1.48 ;
        RECT 3.04 1.24 4.02 1.48 ;
        RECT 3.8 1.48 4.26 1.58 ;
        RECT 3.04 3.56 3.44 4.68 ;
        RECT 3.04 1.08 3.44 1.48 ;
        RECT 3.05 1.08 3.29 4.68 ;
    END
  END AUS
  PIN EIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9552 LAYER ME1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9168 LAYER ME1 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER VI1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME1 ;
      ANTENNAGATEAREA 0.6552 LAYER ME2 ;
      ANTENNAMAXAREACAR 1.457875 LAYER ME1 ;
      ANTENNAMAXAREACAR 1.457875 LAYER ME2 ;
      ANTENNAMAXSIDEAREACAR 5.978022 LAYER ME1 ;
      ANTENNAMAXSIDEAREACAR 5.978022 LAYER ME2 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI1 ;
      ANTENNAMAXCUTCAR 0.119658 LAYER VI2 ;
    PORT
      LAYER VI1 ;
        RECT 1.66 2.02 1.94 2.3 ;
      LAYER ME2 ;
        RECT 1.58 1.94 2.02 2.38 ;
      LAYER ME1 ;
        RECT 1.58 1.94 2.02 2.38 ;
    END
  END EIN0
  PIN vddb
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 5.56 6.48 5.96 ;
    END
  END vddb
  PIN vddd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ME1 ;
        RECT 1.6 3.56 2 5.32 ;
        RECT 4.48 3.56 4.88 5.32 ;
        RECT 0 4.92 6.48 5.32 ;
    END
  END vddd
  PIN gndb
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER ME1 ;
        RECT 0 -0.2 6.48 0.2 ;
    END
  END gndb
  PIN gndd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME1 ;
        RECT 1.6 0.44 2 1.48 ;
        RECT 4.48 0.44 4.88 1.48 ;
        RECT 0 0.44 6.48 0.84 ;
    END
  END gndd
  OBS
    LAYER ME1 ;
      RECT 0.88 1.08 1.28 1.48 ;
      RECT 0.57 2.8 1.17 3.2 ;
      RECT 0.93 1.08 1.17 4.68 ;
      RECT 0.88 3.56 1.28 4.68 ;
      RECT 2.32 1.08 2.72 1.48 ;
      RECT 2.39 2.21 2.79 2.61 ;
      RECT 2.43 1.08 2.67 4.68 ;
      RECT 2.32 3.56 2.72 4.68 ;
      RECT 3.57 2 3.97 2.44 ;
      RECT 3.57 2.2 5.07 2.44 ;
      RECT 4.67 2.2 5.07 2.69 ;
      RECT 5.35 2.38 5.75 2.78 ;
      RECT 3.53 2.8 3.93 3.2 ;
      RECT 5.35 2.38 5.59 3.2 ;
      RECT 3.53 2.96 5.59 3.2 ;
  END
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY filterSize 3 ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY ySnapSpacing 0.01 ;
  PROPERTY xSnapSpacing 0.01 ;
  PROPERTY gridMultiple 1 ;
  PROPERTY gridSpacing 0.72 ;
  PROPERTY stopLevel 32 ;
  PROPERTY startLevel 0 ;
  PROPERTY instLabel "master" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY pathCL "yes" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY instanceDrawingMode "BBox" ;
END UCL_XOR

END LIBRARY
